
library IEEE;
	use IEEE.std_logic_1164.all;
	use IEEE.numeric_std.all;

entity Wrapper_SmallROM is
	port (
		address	: in	std_logic_vector(7 downto 0);
		value	: out	std_logic_vector(7 downto 0)
	);
end entity;

architecture Arch of Wrapper_SmallROM is

	type ROM_t is array (natural range 0 to 255) of std_logic_vector(7 downto 0);
	constant ROM: ROM_t := (
		0 => "11111111",
		1 => "11111110",
		2 => "11111101",
		3 => "11111100",
		4 => "11111011",
		5 => "11111010",
		6 => "11111001",
		7 => "11111000",
		8 => "11110111",
		9 => "11110110",
		10 => "11110101",
		11 => "11110100",
		12 => "11110011",
		13 => "11110010",
		14 => "11110001",
		15 => "11110000",
		16 => "11101111",
		17 => "11101110",
		18 => "11101101",
		19 => "11101100",
		20 => "11101011",
		21 => "11101010",
		22 => "11101001",
		23 => "11101000",
		24 => "11100111",
		25 => "11100110",
		26 => "11100101",
		27 => "11100100",
		28 => "11100011",
		29 => "11100010",
		30 => "11100001",
		31 => "11100000",
		32 => "11011111",
		33 => "11011110",
		34 => "11011101",
		35 => "11011100",
		36 => "11011011",
		37 => "11011010",
		38 => "11011001",
		39 => "11011000",
		40 => "11010111",
		41 => "11010110",
		42 => "11010101",
		43 => "11010100",
		44 => "11010011",
		45 => "11010010",
		46 => "11010001",
		47 => "11010000",
		48 => "11001111",
		49 => "11001110",
		50 => "11001101",
		51 => "11001100",
		52 => "11001011",
		53 => "11001010",
		54 => "11001001",
		55 => "11001000",
		56 => "11000111",
		57 => "11000110",
		58 => "11000101",
		59 => "11000100",
		60 => "11000011",
		61 => "11000010",
		62 => "11000001",
		63 => "11000000",
		64 => "10111111",
		65 => "10111110",
		66 => "10111101",
		67 => "10111100",
		68 => "10111011",
		69 => "10111010",
		70 => "10111001",
		71 => "10111000",
		72 => "10110111",
		73 => "10110110",
		74 => "10110101",
		75 => "10110100",
		76 => "10110011",
		77 => "10110010",
		78 => "10110001",
		79 => "10110000",
		80 => "10101111",
		81 => "10101110",
		82 => "10101101",
		83 => "10101100",
		84 => "10101011",
		85 => "10101010",
		86 => "10101001",
		87 => "10101000",
		88 => "10100111",
		89 => "10100110",
		90 => "10100101",
		91 => "10100100",
		92 => "10100011",
		93 => "10100010",
		94 => "10100001",
		95 => "10100000",
		96 => "10011111",
		97 => "10011110",
		98 => "10011101",
		99 => "10011100",
		100 => "10011011",
		101 => "10011010",
		102 => "10011001",
		103 => "10011000",
		104 => "10010111",
		105 => "10010110",
		106 => "10010101",
		107 => "10010100",
		108 => "10010011",
		109 => "10010010",
		110 => "10010001",
		111 => "10010000",
		112 => "10001111",
		113 => "10001110",
		114 => "10001101",
		115 => "10001100",
		116 => "10001011",
		117 => "10001010",
		118 => "10001001",
		119 => "10001000",
		120 => "10000111",
		121 => "10000110",
		122 => "10000101",
		123 => "10000100",
		124 => "10000011",
		125 => "10000010",
		126 => "10000001",
		127 => "10000000",
		128 => "01111111",
		129 => "01111110",
		130 => "01111101",
		131 => "01111100",
		132 => "01111011",
		133 => "01111010",
		134 => "01111001",
		135 => "01111000",
		136 => "01110111",
		137 => "01110110",
		138 => "01110101",
		139 => "01110100",
		140 => "01110011",
		141 => "01110010",
		142 => "01110001",
		143 => "01110000",
		144 => "01101111",
		145 => "01101110",
		146 => "01101101",
		147 => "01101100",
		148 => "01101011",
		149 => "01101010",
		150 => "01101001",
		151 => "01101000",
		152 => "01100111",
		153 => "01100110",
		154 => "01100101",
		155 => "01100100",
		156 => "01100011",
		157 => "01100010",
		158 => "01100001",
		159 => "01100000",
		160 => "01011111",
		161 => "01011110",
		162 => "01011101",
		163 => "01011100",
		164 => "01011011",
		165 => "01011010",
		166 => "01011001",
		167 => "01011000",
		168 => "01010111",
		169 => "01010110",
		170 => "01010101",
		171 => "01010100",
		172 => "01010011",
		173 => "01010010",
		174 => "01010001",
		175 => "01010000",
		176 => "01001111",
		177 => "01001110",
		178 => "01001101",
		179 => "01001100",
		180 => "01001011",
		181 => "01001010",
		182 => "01001001",
		183 => "01001000",
		184 => "01000111",
		185 => "01000110",
		186 => "01000101",
		187 => "01000100",
		188 => "01000011",
		189 => "01000010",
		190 => "01000001",
		191 => "01000000",
		192 => "00111111",
		193 => "00111110",
		194 => "00111101",
		195 => "00111100",
		196 => "00111011",
		197 => "00111010",
		198 => "00111001",
		199 => "00111000",
		200 => "00110111",
		201 => "00110110",
		202 => "00110101",
		203 => "00110100",
		204 => "00110011",
		205 => "00110010",
		206 => "00110001",
		207 => "00110000",
		208 => "00101111",
		209 => "00101110",
		210 => "00101101",
		211 => "00101100",
		212 => "00101011",
		213 => "00101010",
		214 => "00101001",
		215 => "00101000",
		216 => "00100111",
		217 => "00100110",
		218 => "00100101",
		219 => "00100100",
		220 => "00100011",
		221 => "00100010",
		222 => "00100001",
		223 => "00100000",
		224 => "00011111",
		225 => "00011110",
		226 => "00011101",
		227 => "00011100",
		228 => "00011011",
		229 => "00011010",
		230 => "00011001",
		231 => "00011000",
		232 => "00010111",
		233 => "00010110",
		234 => "00010101",
		235 => "00010100",
		236 => "00010011",
		237 => "00010010",
		238 => "00010001",
		239 => "00010000",
		240 => "00001111",
		241 => "00001110",
		242 => "00001101",
		243 => "00001100",
		244 => "00001011",
		245 => "00001010",
		246 => "00001001",
		247 => "00001000",
		248 => "00000111",
		249 => "00000110",
		250 => "00000101",
		251 => "00000100",
		252 => "00000011",
		253 => "00000010",
		254 => "00000001",
		255 => "00000000"
	);

begin

	value <= ROM( to_integer( unsigned(address) ) );

end architecture;
