
library IEEE;
	use IEEE.std_logic_1164.all;
	use IEEE.numeric_std.all;

entity ROM is
	port (
		address	: in	std_logic_vector(13 downto 0);
		value	: out	std_logic_vector(7 downto 0)
	);
end entity;

architecture Arch of ROM is

	type ROM_t is array (natural range 0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM: ROM_t := (
		0 => "11111111",
		1 => "11111111",
		2 => "11111111",
		3 => "11111111",
		4 => "11111111",
		5 => "11111111",
		6 => "11111111",
		7 => "11111111",
		8 => "11111111",
		9 => "11111111",
		10 => "11111111",
		11 => "11111111",
		12 => "11111111",
		13 => "11111111",
		14 => "11111111",
		15 => "11111111",
		16 => "11111111",
		17 => "11111111",
		18 => "11111111",
		19 => "11111111",
		20 => "11111111",
		21 => "11111111",
		22 => "11111111",
		23 => "11111111",
		24 => "11111111",
		25 => "11111111",
		26 => "11111111",
		27 => "11111111",
		28 => "11111111",
		29 => "11111111",
		30 => "11111111",
		31 => "11111111",
		32 => "11111111",
		33 => "11111111",
		34 => "11111111",
		35 => "11111111",
		36 => "11111111",
		37 => "11111111",
		38 => "11111111",
		39 => "11111111",
		40 => "11111111",
		41 => "11111111",
		42 => "11111111",
		43 => "11111111",
		44 => "11111111",
		45 => "11111111",
		46 => "11111111",
		47 => "11111111",
		48 => "11111111",
		49 => "11111111",
		50 => "11111111",
		51 => "11111111",
		52 => "11111111",
		53 => "11111111",
		54 => "11111111",
		55 => "11111111",
		56 => "11111111",
		57 => "11111111",
		58 => "11111111",
		59 => "11111111",
		60 => "11111111",
		61 => "11111111",
		62 => "11111111",
		63 => "11111111",
		64 => "11111111",
		65 => "11111111",
		66 => "11111111",
		67 => "11111111",
		68 => "11111111",
		69 => "11111111",
		70 => "11111111",
		71 => "11111111",
		72 => "11111111",
		73 => "11111111",
		74 => "11111111",
		75 => "11111111",
		76 => "11111111",
		77 => "11111111",
		78 => "11111111",
		79 => "11111111",
		80 => "11111111",
		81 => "11111111",
		82 => "11111111",
		83 => "11111111",
		84 => "11111111",
		85 => "11111111",
		86 => "11111111",
		87 => "11111111",
		88 => "11111111",
		89 => "11111111",
		90 => "11111111",
		91 => "11111111",
		92 => "11111111",
		93 => "11111111",
		94 => "11111111",
		95 => "11111111",
		96 => "11111111",
		97 => "11111111",
		98 => "11111111",
		99 => "11111111",
		100 => "11111111",
		101 => "11111111",
		102 => "11111111",
		103 => "11111111",
		104 => "11111111",
		105 => "11111111",
		106 => "11111111",
		107 => "11111111",
		108 => "11111111",
		109 => "11111111",
		110 => "11111111",
		111 => "11111111",
		112 => "11111111",
		113 => "11111111",
		114 => "11111111",
		115 => "11111111",
		116 => "11111111",
		117 => "11111111",
		118 => "11111111",
		119 => "11111111",
		120 => "11111111",
		121 => "11111111",
		122 => "11111111",
		123 => "11111111",
		124 => "11111111",
		125 => "11111111",
		126 => "11111111",
		127 => "11111111",
		128 => "11111111",
		129 => "11111111",
		130 => "11111111",
		131 => "11111111",
		132 => "11111111",
		133 => "11111111",
		134 => "11111111",
		135 => "11111111",
		136 => "11111111",
		137 => "11111111",
		138 => "11111111",
		139 => "11111111",
		140 => "11111111",
		141 => "11111111",
		142 => "11111111",
		143 => "11111111",
		144 => "11111111",
		145 => "11111111",
		146 => "11111111",
		147 => "11111111",
		148 => "11111111",
		149 => "11111111",
		150 => "11111111",
		151 => "11111111",
		152 => "11111111",
		153 => "11111111",
		154 => "11111111",
		155 => "11111111",
		156 => "11111111",
		157 => "11111111",
		158 => "11111111",
		159 => "11111111",
		160 => "11111111",
		161 => "11111111",
		162 => "11111111",
		163 => "11111111",
		164 => "11111111",
		165 => "11111111",
		166 => "11111111",
		167 => "11111111",
		168 => "11111111",
		169 => "11111111",
		170 => "11111111",
		171 => "11111111",
		172 => "11111111",
		173 => "11111111",
		174 => "11111111",
		175 => "11111111",
		176 => "11111111",
		177 => "11111111",
		178 => "11111111",
		179 => "11111111",
		180 => "11111111",
		181 => "11111111",
		182 => "11111111",
		183 => "11111111",
		184 => "11111111",
		185 => "11111111",
		186 => "11111111",
		187 => "11111111",
		188 => "11111111",
		189 => "11111111",
		190 => "11111111",
		191 => "11111111",
		192 => "11111111",
		193 => "11111111",
		194 => "11111111",
		195 => "11111111",
		196 => "11111111",
		197 => "11111111",
		198 => "11111111",
		199 => "11111111",
		200 => "11111111",
		201 => "11111111",
		202 => "11111111",
		203 => "11111111",
		204 => "11111111",
		205 => "11111111",
		206 => "11111111",
		207 => "11111111",
		208 => "11111111",
		209 => "11111111",
		210 => "11111111",
		211 => "11111111",
		212 => "11111111",
		213 => "11111111",
		214 => "11111111",
		215 => "11111111",
		216 => "11111111",
		217 => "11111111",
		218 => "11111111",
		219 => "11111111",
		220 => "11111111",
		221 => "11111111",
		222 => "11111111",
		223 => "11111111",
		224 => "11111111",
		225 => "11111111",
		226 => "11111111",
		227 => "11111111",
		228 => "11111111",
		229 => "11111111",
		230 => "11111111",
		231 => "11111111",
		232 => "11111111",
		233 => "11111111",
		234 => "11111111",
		235 => "11111111",
		236 => "11111111",
		237 => "11111111",
		238 => "11111111",
		239 => "11111111",
		240 => "11111111",
		241 => "11111111",
		242 => "11111111",
		243 => "11111111",
		244 => "11111111",
		245 => "11111111",
		246 => "11111111",
		247 => "11111111",
		248 => "11111111",
		249 => "11111111",
		250 => "11111111",
		251 => "11111111",
		252 => "11111111",
		253 => "11111111",
		254 => "11111111",
		255 => "11111111",
		256 => "11111111",
		257 => "11111111",
		258 => "11111111",
		259 => "11111111",
		260 => "11111111",
		261 => "11111111",
		262 => "11111111",
		263 => "11111111",
		264 => "11111111",
		265 => "11111111",
		266 => "11111111",
		267 => "11111111",
		268 => "11111111",
		269 => "11111111",
		270 => "11111111",
		271 => "11111111",
		272 => "11111111",
		273 => "11111111",
		274 => "11111111",
		275 => "11111111",
		276 => "11111111",
		277 => "11111111",
		278 => "11111111",
		279 => "11111111",
		280 => "11111111",
		281 => "11111111",
		282 => "11111111",
		283 => "11111111",
		284 => "11111111",
		285 => "11111111",
		286 => "11111111",
		287 => "11111111",
		288 => "11111111",
		289 => "11111111",
		290 => "11111111",
		291 => "11111111",
		292 => "11111111",
		293 => "11111111",
		294 => "11111111",
		295 => "11111111",
		296 => "11111111",
		297 => "11111111",
		298 => "11111111",
		299 => "11111111",
		300 => "11111111",
		301 => "11111111",
		302 => "11111111",
		303 => "11111111",
		304 => "11111111",
		305 => "11111111",
		306 => "11111111",
		307 => "11111111",
		308 => "11111111",
		309 => "11111111",
		310 => "11111111",
		311 => "11111111",
		312 => "11111111",
		313 => "11111111",
		314 => "11111111",
		315 => "11111111",
		316 => "11111111",
		317 => "11111111",
		318 => "11111111",
		319 => "11111111",
		320 => "11111111",
		321 => "11111111",
		322 => "11111111",
		323 => "11111111",
		324 => "11111111",
		325 => "11111111",
		326 => "11111111",
		327 => "11111111",
		328 => "11111111",
		329 => "11111111",
		330 => "11111111",
		331 => "11111111",
		332 => "11111111",
		333 => "11111111",
		334 => "11111111",
		335 => "11111111",
		336 => "11111111",
		337 => "11111111",
		338 => "11111111",
		339 => "11111111",
		340 => "11111111",
		341 => "11111111",
		342 => "11111111",
		343 => "11111111",
		344 => "11111111",
		345 => "11111111",
		346 => "11111111",
		347 => "11111111",
		348 => "11111111",
		349 => "11111111",
		350 => "11111111",
		351 => "11111111",
		352 => "11111111",
		353 => "11111111",
		354 => "11111111",
		355 => "11111111",
		356 => "11111111",
		357 => "11111111",
		358 => "11111111",
		359 => "11111111",
		360 => "11111111",
		361 => "11111111",
		362 => "11111111",
		363 => "11111111",
		364 => "11111111",
		365 => "11111111",
		366 => "11111111",
		367 => "11111111",
		368 => "11111111",
		369 => "11111111",
		370 => "11111111",
		371 => "11111111",
		372 => "11111111",
		373 => "11111111",
		374 => "11111111",
		375 => "11111111",
		376 => "11111111",
		377 => "11111111",
		378 => "11111111",
		379 => "11111111",
		380 => "11111111",
		381 => "11111111",
		382 => "11111111",
		383 => "11111111",
		384 => "11111111",
		385 => "11111111",
		386 => "11111111",
		387 => "11111111",
		388 => "11111111",
		389 => "11111111",
		390 => "11111111",
		391 => "11111111",
		392 => "11111111",
		393 => "11111111",
		394 => "11111111",
		395 => "11111111",
		396 => "11111111",
		397 => "11111111",
		398 => "11111111",
		399 => "11111111",
		400 => "11111111",
		401 => "11111111",
		402 => "11111111",
		403 => "11111111",
		404 => "11111111",
		405 => "11111111",
		406 => "11111111",
		407 => "11111111",
		408 => "11111111",
		409 => "11111111",
		410 => "11111111",
		411 => "11111111",
		412 => "11111111",
		413 => "11111111",
		414 => "11111111",
		415 => "11111111",
		416 => "11111111",
		417 => "11111111",
		418 => "11111111",
		419 => "11111111",
		420 => "11111111",
		421 => "11111111",
		422 => "11111111",
		423 => "11111111",
		424 => "11111111",
		425 => "11111111",
		426 => "11111111",
		427 => "11111111",
		428 => "11111111",
		429 => "11111111",
		430 => "11111111",
		431 => "11111111",
		432 => "11111111",
		433 => "11111111",
		434 => "11111111",
		435 => "11111111",
		436 => "11111111",
		437 => "11111111",
		438 => "11111111",
		439 => "11111111",
		440 => "11111111",
		441 => "11111111",
		442 => "11111111",
		443 => "11111111",
		444 => "11111111",
		445 => "11111111",
		446 => "11111111",
		447 => "11111111",
		448 => "11111111",
		449 => "11111111",
		450 => "11111111",
		451 => "11111111",
		452 => "11111111",
		453 => "11111111",
		454 => "11111111",
		455 => "11111111",
		456 => "11111111",
		457 => "11111111",
		458 => "11111111",
		459 => "11111111",
		460 => "11111111",
		461 => "11111111",
		462 => "11111111",
		463 => "11111111",
		464 => "11111111",
		465 => "11111111",
		466 => "11111111",
		467 => "11111111",
		468 => "11111111",
		469 => "11111111",
		470 => "11111111",
		471 => "11111111",
		472 => "11111111",
		473 => "11111111",
		474 => "11111111",
		475 => "11111111",
		476 => "11111111",
		477 => "11111111",
		478 => "11111111",
		479 => "11111111",
		480 => "11111111",
		481 => "11111111",
		482 => "11111111",
		483 => "11111111",
		484 => "11111111",
		485 => "11111111",
		486 => "11111111",
		487 => "11111111",
		488 => "11111111",
		489 => "11111111",
		490 => "11111111",
		491 => "11111111",
		492 => "11111111",
		493 => "11111111",
		494 => "11111111",
		495 => "11111111",
		496 => "11111111",
		497 => "11111111",
		498 => "11111111",
		499 => "11111111",
		500 => "11111111",
		501 => "11111111",
		502 => "11111111",
		503 => "11111111",
		504 => "11111111",
		505 => "11111111",
		506 => "11111111",
		507 => "11111111",
		508 => "11111111",
		509 => "11111111",
		510 => "11111111",
		511 => "11111111",
		512 => "11111111",
		513 => "11111111",
		514 => "11111111",
		515 => "11111111",
		516 => "11111111",
		517 => "11111111",
		518 => "11111111",
		519 => "11111111",
		520 => "11111111",
		521 => "11111111",
		522 => "11111111",
		523 => "11111111",
		524 => "11111111",
		525 => "11111111",
		526 => "11111111",
		527 => "11111111",
		528 => "11111111",
		529 => "11111111",
		530 => "11111111",
		531 => "11111111",
		532 => "11111111",
		533 => "11111111",
		534 => "11111111",
		535 => "11111111",
		536 => "11111111",
		537 => "11111111",
		538 => "11111111",
		539 => "11111111",
		540 => "11111111",
		541 => "11111111",
		542 => "11111111",
		543 => "11111111",
		544 => "11111111",
		545 => "11111111",
		546 => "11111111",
		547 => "11111111",
		548 => "11111111",
		549 => "11111111",
		550 => "11111111",
		551 => "11111111",
		552 => "11111111",
		553 => "11111111",
		554 => "11111111",
		555 => "11111111",
		556 => "11111111",
		557 => "11111111",
		558 => "11111111",
		559 => "11111111",
		560 => "11111111",
		561 => "11111111",
		562 => "11111111",
		563 => "11111111",
		564 => "11111111",
		565 => "11111111",
		566 => "11111111",
		567 => "11111111",
		568 => "11100010",
		569 => "11010001",
		570 => "10101110",
		571 => "10100011",
		572 => "01111100",
		573 => "01110101",
		574 => "01010011",
		575 => "11111111",
		576 => "11111111",
		577 => "11111111",
		578 => "11111111",
		579 => "11111111",
		580 => "11111111",
		581 => "11111111",
		582 => "11111111",
		583 => "11111111",
		584 => "11111111",
		585 => "11111111",
		586 => "11111111",
		587 => "11111111",
		588 => "11111111",
		589 => "11111111",
		590 => "11111111",
		591 => "11111111",
		592 => "11111111",
		593 => "11111111",
		594 => "11111111",
		595 => "11111111",
		596 => "11111111",
		597 => "11111111",
		598 => "11111111",
		599 => "11111111",
		600 => "11111111",
		601 => "11111111",
		602 => "11111111",
		603 => "11111111",
		604 => "11111111",
		605 => "11111111",
		606 => "11111111",
		607 => "11111111",
		608 => "11111111",
		609 => "11111111",
		610 => "11111111",
		611 => "11111111",
		612 => "11111111",
		613 => "11111111",
		614 => "11111111",
		615 => "11111111",
		616 => "11111111",
		617 => "11111111",
		618 => "11111111",
		619 => "11111111",
		620 => "11111111",
		621 => "11111111",
		622 => "11111111",
		623 => "11111111",
		624 => "11111111",
		625 => "11111111",
		626 => "11111111",
		627 => "11111111",
		628 => "11111111",
		629 => "11111111",
		630 => "11111111",
		631 => "11111111",
		632 => "11111111",
		633 => "11111111",
		634 => "11111111",
		635 => "11111111",
		636 => "11111111",
		637 => "11111111",
		638 => "11111111",
		639 => "11111111",
		640 => "11111111",
		641 => "11111111",
		642 => "11111111",
		643 => "11111111",
		644 => "11111111",
		645 => "11111111",
		646 => "11111111",
		647 => "11111111",
		648 => "11111111",
		649 => "11111111",
		650 => "11111111",
		651 => "11111111",
		652 => "11111111",
		653 => "11111111",
		654 => "11111111",
		655 => "11111111",
		656 => "11111111",
		657 => "11111111",
		658 => "11111111",
		659 => "11111111",
		660 => "11111111",
		661 => "11111111",
		662 => "11111111",
		663 => "11111111",
		664 => "11111111",
		665 => "11111111",
		666 => "11111111",
		667 => "11111111",
		668 => "11111111",
		669 => "11111111",
		670 => "11111111",
		671 => "11111111",
		672 => "11111111",
		673 => "11111111",
		674 => "11111111",
		675 => "11111111",
		676 => "11111111",
		677 => "11111111",
		678 => "11111111",
		679 => "11111111",
		680 => "11111111",
		681 => "11111111",
		682 => "11111111",
		683 => "11111111",
		684 => "11111111",
		685 => "11111111",
		686 => "11111111",
		687 => "11111111",
		688 => "11111111",
		689 => "11111111",
		690 => "11111111",
		691 => "11111111",
		692 => "11111111",
		693 => "11111111",
		694 => "11111111",
		695 => "01110101",
		696 => "01000111",
		697 => "01011110",
		698 => "11000101",
		699 => "11010001",
		700 => "11111111",
		701 => "11010111",
		702 => "01000111",
		703 => "11110011",
		704 => "11111111",
		705 => "11111111",
		706 => "11111111",
		707 => "11111111",
		708 => "11111111",
		709 => "11111111",
		710 => "11111111",
		711 => "11111111",
		712 => "11111111",
		713 => "11111111",
		714 => "11010001",
		715 => "01110101",
		716 => "10100011",
		717 => "11010111",
		718 => "11111111",
		719 => "11111111",
		720 => "11111111",
		721 => "11111111",
		722 => "11111111",
		723 => "11111111",
		724 => "11111111",
		725 => "11111111",
		726 => "11111111",
		727 => "11111111",
		728 => "11111111",
		729 => "11111111",
		730 => "11111111",
		731 => "11111111",
		732 => "11111111",
		733 => "11111111",
		734 => "11111111",
		735 => "11111111",
		736 => "11111111",
		737 => "11111111",
		738 => "11111111",
		739 => "11111111",
		740 => "11111111",
		741 => "11111111",
		742 => "11111111",
		743 => "11111111",
		744 => "11111111",
		745 => "11111111",
		746 => "11111111",
		747 => "11111111",
		748 => "11111111",
		749 => "11111111",
		750 => "11111111",
		751 => "11111111",
		752 => "11111111",
		753 => "11111111",
		754 => "11111111",
		755 => "11111111",
		756 => "11111111",
		757 => "11111111",
		758 => "11111111",
		759 => "11111111",
		760 => "11111111",
		761 => "11111111",
		762 => "11111111",
		763 => "11111111",
		764 => "11111111",
		765 => "11111111",
		766 => "11111111",
		767 => "11111111",
		768 => "11111111",
		769 => "11111111",
		770 => "11111111",
		771 => "11111111",
		772 => "11111111",
		773 => "11111111",
		774 => "11111111",
		775 => "11111111",
		776 => "11111111",
		777 => "11111111",
		778 => "11111111",
		779 => "11111111",
		780 => "11111111",
		781 => "11111111",
		782 => "11111111",
		783 => "11111111",
		784 => "11111111",
		785 => "11111111",
		786 => "11111111",
		787 => "11111111",
		788 => "11111111",
		789 => "11111111",
		790 => "11111111",
		791 => "11111111",
		792 => "11111111",
		793 => "11111111",
		794 => "11111111",
		795 => "11111111",
		796 => "11111111",
		797 => "11111111",
		798 => "11111111",
		799 => "11111111",
		800 => "11111111",
		801 => "11111111",
		802 => "11111111",
		803 => "11111111",
		804 => "11111111",
		805 => "11111111",
		806 => "11111111",
		807 => "11111111",
		808 => "11111111",
		809 => "11111111",
		810 => "11111111",
		811 => "11111111",
		812 => "11111111",
		813 => "11111111",
		814 => "11111111",
		815 => "11111111",
		816 => "11111111",
		817 => "11111111",
		818 => "11111111",
		819 => "11111111",
		820 => "11111111",
		821 => "11111111",
		822 => "11101000",
		823 => "01110101",
		824 => "01011001",
		825 => "01011001",
		826 => "11111111",
		827 => "11111111",
		828 => "11111111",
		829 => "11111111",
		830 => "10011110",
		831 => "11100010",
		832 => "11111111",
		833 => "11111111",
		834 => "11111111",
		835 => "11111111",
		836 => "11111111",
		837 => "11111111",
		838 => "11111111",
		839 => "11111111",
		840 => "11111111",
		841 => "11111111",
		842 => "11111111",
		843 => "11010001",
		844 => "01000111",
		845 => "01010011",
		846 => "01011110",
		847 => "10000111",
		848 => "10111010",
		849 => "11111001",
		850 => "11111111",
		851 => "11111111",
		852 => "11111111",
		853 => "11111111",
		854 => "11111111",
		855 => "11111111",
		856 => "11111111",
		857 => "11111111",
		858 => "11111111",
		859 => "11111111",
		860 => "11111111",
		861 => "11111111",
		862 => "11111111",
		863 => "11111111",
		864 => "11111111",
		865 => "11111111",
		866 => "11111111",
		867 => "11111111",
		868 => "11111111",
		869 => "11111111",
		870 => "11111111",
		871 => "11111111",
		872 => "11111111",
		873 => "11111111",
		874 => "11111111",
		875 => "11111111",
		876 => "11111111",
		877 => "11111111",
		878 => "11111111",
		879 => "11111111",
		880 => "11111111",
		881 => "11111111",
		882 => "11111111",
		883 => "11111111",
		884 => "11111111",
		885 => "11111111",
		886 => "11111111",
		887 => "11111111",
		888 => "11111111",
		889 => "11111111",
		890 => "11111111",
		891 => "11111111",
		892 => "11111111",
		893 => "11111111",
		894 => "11111111",
		895 => "11111111",
		896 => "11111111",
		897 => "11111111",
		898 => "11111111",
		899 => "11111111",
		900 => "11111111",
		901 => "11111111",
		902 => "11111111",
		903 => "11111111",
		904 => "11111111",
		905 => "11111111",
		906 => "11111111",
		907 => "11111111",
		908 => "11111111",
		909 => "11111111",
		910 => "11111111",
		911 => "11111111",
		912 => "11111111",
		913 => "11111111",
		914 => "11111111",
		915 => "11111111",
		916 => "11111111",
		917 => "11111111",
		918 => "11111111",
		919 => "11111111",
		920 => "11111111",
		921 => "11111111",
		922 => "11111111",
		923 => "11111111",
		924 => "11111111",
		925 => "11111111",
		926 => "11111111",
		927 => "11111111",
		928 => "11111111",
		929 => "11111111",
		930 => "11111111",
		931 => "11111111",
		932 => "11111111",
		933 => "11111111",
		934 => "11111111",
		935 => "11111111",
		936 => "11111111",
		937 => "11111111",
		938 => "11111111",
		939 => "11101110",
		940 => "10011110",
		941 => "11111111",
		942 => "11111111",
		943 => "11111111",
		944 => "11111111",
		945 => "11111111",
		946 => "11111111",
		947 => "11111111",
		948 => "11111111",
		949 => "11111111",
		950 => "10100011",
		951 => "10110100",
		952 => "01110000",
		953 => "01000111",
		954 => "11111001",
		955 => "11111111",
		956 => "11111111",
		957 => "11111111",
		958 => "11111111",
		959 => "11111111",
		960 => "11111111",
		961 => "11111111",
		962 => "11111111",
		963 => "11111111",
		964 => "11111111",
		965 => "11111111",
		966 => "11111111",
		967 => "11111111",
		968 => "11111111",
		969 => "11111111",
		970 => "11111111",
		971 => "10111010",
		972 => "01000111",
		973 => "10011110",
		974 => "11111111",
		975 => "11011100",
		976 => "10001100",
		977 => "01010011",
		978 => "10100011",
		979 => "11111111",
		980 => "11111111",
		981 => "11111111",
		982 => "11111111",
		983 => "11111111",
		984 => "11111111",
		985 => "11111111",
		986 => "11111111",
		987 => "11111111",
		988 => "11111111",
		989 => "11111111",
		990 => "11111111",
		991 => "11111111",
		992 => "11111111",
		993 => "11111111",
		994 => "11111111",
		995 => "11111111",
		996 => "11111111",
		997 => "11111111",
		998 => "11111111",
		999 => "11111111",
		1000 => "11111111",
		1001 => "11111111",
		1002 => "11111111",
		1003 => "11111111",
		1004 => "11111111",
		1005 => "11111111",
		1006 => "11111111",
		1007 => "11111111",
		1008 => "11111111",
		1009 => "11111111",
		1010 => "11111111",
		1011 => "11111111",
		1012 => "11111111",
		1013 => "11111111",
		1014 => "11111111",
		1015 => "11111111",
		1016 => "11111111",
		1017 => "11111111",
		1018 => "11111111",
		1019 => "11111111",
		1020 => "11111111",
		1021 => "11111111",
		1022 => "11111111",
		1023 => "11111111",
		1024 => "11111111",
		1025 => "11111111",
		1026 => "11111111",
		1027 => "11111111",
		1028 => "11111111",
		1029 => "11111111",
		1030 => "11111111",
		1031 => "11111111",
		1032 => "11111111",
		1033 => "11111111",
		1034 => "11111111",
		1035 => "11111111",
		1036 => "11111111",
		1037 => "11111111",
		1038 => "11111111",
		1039 => "11111111",
		1040 => "11111111",
		1041 => "11111111",
		1042 => "11111111",
		1043 => "11111111",
		1044 => "11111111",
		1045 => "11111111",
		1046 => "11111111",
		1047 => "11111111",
		1048 => "11111111",
		1049 => "11111111",
		1050 => "11111111",
		1051 => "11111111",
		1052 => "11111111",
		1053 => "11111111",
		1054 => "11111111",
		1055 => "11111111",
		1056 => "11111111",
		1057 => "11111111",
		1058 => "11111111",
		1059 => "11111111",
		1060 => "11111111",
		1061 => "11111111",
		1062 => "11111111",
		1063 => "11111111",
		1064 => "11111111",
		1065 => "11101110",
		1066 => "10011000",
		1067 => "01001101",
		1068 => "10111010",
		1069 => "11111111",
		1070 => "11111111",
		1071 => "11111111",
		1072 => "11111111",
		1073 => "11111111",
		1074 => "11111111",
		1075 => "11111111",
		1076 => "11111111",
		1077 => "11111111",
		1078 => "01011110",
		1079 => "11101110",
		1080 => "10000111",
		1081 => "01000111",
		1082 => "11100010",
		1083 => "11111111",
		1084 => "11111111",
		1085 => "11101110",
		1086 => "10111010",
		1087 => "11111111",
		1088 => "11111111",
		1089 => "11111111",
		1090 => "11111111",
		1091 => "11111111",
		1092 => "11111111",
		1093 => "11111111",
		1094 => "11111111",
		1095 => "11111111",
		1096 => "11111111",
		1097 => "11111111",
		1098 => "11111111",
		1099 => "10001100",
		1100 => "01000111",
		1101 => "11010001",
		1102 => "11111111",
		1103 => "11111111",
		1104 => "11111111",
		1105 => "11100010",
		1106 => "01001101",
		1107 => "10011000",
		1108 => "11111111",
		1109 => "11111111",
		1110 => "11111111",
		1111 => "11111111",
		1112 => "11111111",
		1113 => "11111111",
		1114 => "11111111",
		1115 => "11111111",
		1116 => "11111111",
		1117 => "11111111",
		1118 => "11111111",
		1119 => "11111111",
		1120 => "11111111",
		1121 => "11111111",
		1122 => "11111111",
		1123 => "11111111",
		1124 => "11111111",
		1125 => "11111111",
		1126 => "11111111",
		1127 => "11111111",
		1128 => "11111111",
		1129 => "11111111",
		1130 => "11111111",
		1131 => "11111111",
		1132 => "11111111",
		1133 => "11111111",
		1134 => "11111111",
		1135 => "11111111",
		1136 => "11111111",
		1137 => "11111111",
		1138 => "11111111",
		1139 => "11111111",
		1140 => "11111111",
		1141 => "11111111",
		1142 => "11111111",
		1143 => "11111111",
		1144 => "11111111",
		1145 => "11111111",
		1146 => "11111111",
		1147 => "11111111",
		1148 => "11111111",
		1149 => "11111111",
		1150 => "11111111",
		1151 => "11111111",
		1152 => "11111111",
		1153 => "11111111",
		1154 => "11111111",
		1155 => "11111111",
		1156 => "11111111",
		1157 => "11111111",
		1158 => "11111111",
		1159 => "11111111",
		1160 => "11111111",
		1161 => "11111111",
		1162 => "11111111",
		1163 => "11111111",
		1164 => "11111111",
		1165 => "11111111",
		1166 => "11111111",
		1167 => "11111111",
		1168 => "11111111",
		1169 => "11111111",
		1170 => "11111111",
		1171 => "11111111",
		1172 => "11111111",
		1173 => "11111111",
		1174 => "11111111",
		1175 => "11111111",
		1176 => "11111111",
		1177 => "11111111",
		1178 => "11111111",
		1179 => "11111111",
		1180 => "11111111",
		1181 => "11111111",
		1182 => "11111111",
		1183 => "11111111",
		1184 => "11111111",
		1185 => "11111111",
		1186 => "11111111",
		1187 => "11111111",
		1188 => "11111111",
		1189 => "11111111",
		1190 => "11111111",
		1191 => "11111111",
		1192 => "11111111",
		1193 => "11000000",
		1194 => "01000111",
		1195 => "01001101",
		1196 => "11101110",
		1197 => "11111111",
		1198 => "11111111",
		1199 => "11111111",
		1200 => "11111111",
		1201 => "11111111",
		1202 => "11111111",
		1203 => "11111111",
		1204 => "11111111",
		1205 => "11111111",
		1206 => "01110101",
		1207 => "11111111",
		1208 => "10100011",
		1209 => "01000111",
		1210 => "11001011",
		1211 => "11111111",
		1212 => "11111111",
		1213 => "11000000",
		1214 => "10000111",
		1215 => "11111111",
		1216 => "11111111",
		1217 => "11111111",
		1218 => "11111111",
		1219 => "11111111",
		1220 => "11111111",
		1221 => "11111111",
		1222 => "11111111",
		1223 => "11111111",
		1224 => "11111111",
		1225 => "11111111",
		1226 => "11111111",
		1227 => "01010011",
		1228 => "01010011",
		1229 => "11111111",
		1230 => "11111111",
		1231 => "11111111",
		1232 => "11111111",
		1233 => "11111111",
		1234 => "10101110",
		1235 => "01000111",
		1236 => "11010001",
		1237 => "11111111",
		1238 => "11111111",
		1239 => "11111111",
		1240 => "11111111",
		1241 => "11111111",
		1242 => "11111111",
		1243 => "11111111",
		1244 => "11111111",
		1245 => "11111111",
		1246 => "11111111",
		1247 => "11111111",
		1248 => "11111111",
		1249 => "11111111",
		1250 => "11111111",
		1251 => "11111111",
		1252 => "11111111",
		1253 => "11111111",
		1254 => "11111111",
		1255 => "11111111",
		1256 => "11111111",
		1257 => "11111111",
		1258 => "11111111",
		1259 => "11111111",
		1260 => "11111111",
		1261 => "11111111",
		1262 => "11111111",
		1263 => "11111111",
		1264 => "11111111",
		1265 => "11111111",
		1266 => "11111111",
		1267 => "11111111",
		1268 => "11111111",
		1269 => "11111111",
		1270 => "11111111",
		1271 => "11111111",
		1272 => "11111111",
		1273 => "11111111",
		1274 => "11111111",
		1275 => "11111111",
		1276 => "11111111",
		1277 => "11111111",
		1278 => "11111111",
		1279 => "11111111",
		1280 => "11111111",
		1281 => "11111111",
		1282 => "11111111",
		1283 => "11111111",
		1284 => "11111111",
		1285 => "11111111",
		1286 => "11111111",
		1287 => "11111111",
		1288 => "11111111",
		1289 => "11111111",
		1290 => "11111111",
		1291 => "11111111",
		1292 => "11111111",
		1293 => "11111111",
		1294 => "11111111",
		1295 => "11111111",
		1296 => "11111111",
		1297 => "11111111",
		1298 => "11111111",
		1299 => "11111111",
		1300 => "11111111",
		1301 => "11111111",
		1302 => "11111111",
		1303 => "11111111",
		1304 => "11111111",
		1305 => "11111111",
		1306 => "11111111",
		1307 => "11111111",
		1308 => "11111111",
		1309 => "11111111",
		1310 => "11111111",
		1311 => "11111111",
		1312 => "11111111",
		1313 => "11111111",
		1314 => "11111111",
		1315 => "11111111",
		1316 => "11111111",
		1317 => "11111111",
		1318 => "11111111",
		1319 => "11111111",
		1320 => "11111111",
		1321 => "11010001",
		1322 => "01001101",
		1323 => "01000111",
		1324 => "10011000",
		1325 => "11111111",
		1326 => "11111111",
		1327 => "11111111",
		1328 => "11111111",
		1329 => "11111111",
		1330 => "11111111",
		1331 => "11111111",
		1332 => "11111111",
		1333 => "11111111",
		1334 => "10110100",
		1335 => "11111111",
		1336 => "10111010",
		1337 => "01000111",
		1338 => "10000001",
		1339 => "10100011",
		1340 => "01110101",
		1341 => "01011110",
		1342 => "01101010",
		1343 => "11111111",
		1344 => "11111111",
		1345 => "11111111",
		1346 => "11111111",
		1347 => "11111111",
		1348 => "11111111",
		1349 => "11111111",
		1350 => "11111111",
		1351 => "11111111",
		1352 => "11111111",
		1353 => "11111111",
		1354 => "11010001",
		1355 => "01000111",
		1356 => "10001100",
		1357 => "11111111",
		1358 => "11111111",
		1359 => "11111111",
		1360 => "11111111",
		1361 => "11111111",
		1362 => "11101110",
		1363 => "01000111",
		1364 => "10010011",
		1365 => "11111111",
		1366 => "11111111",
		1367 => "11111111",
		1368 => "11111111",
		1369 => "11111111",
		1370 => "10101001",
		1371 => "11011100",
		1372 => "11111111",
		1373 => "11111111",
		1374 => "11111111",
		1375 => "11111111",
		1376 => "11111111",
		1377 => "11111111",
		1378 => "11111111",
		1379 => "11111111",
		1380 => "11111111",
		1381 => "11111111",
		1382 => "11111111",
		1383 => "11111111",
		1384 => "11111111",
		1385 => "11111111",
		1386 => "11111111",
		1387 => "11111111",
		1388 => "11111111",
		1389 => "11111111",
		1390 => "11111111",
		1391 => "11111111",
		1392 => "11111111",
		1393 => "11111111",
		1394 => "11111111",
		1395 => "11111111",
		1396 => "11111111",
		1397 => "11111111",
		1398 => "11111111",
		1399 => "11111111",
		1400 => "11111111",
		1401 => "11111111",
		1402 => "11111111",
		1403 => "11111111",
		1404 => "11111111",
		1405 => "11111111",
		1406 => "11111111",
		1407 => "11111111",
		1408 => "11111111",
		1409 => "11111111",
		1410 => "11111111",
		1411 => "11111111",
		1412 => "11111111",
		1413 => "11111111",
		1414 => "11111111",
		1415 => "11111111",
		1416 => "11111111",
		1417 => "11111111",
		1418 => "11111111",
		1419 => "11111111",
		1420 => "11111111",
		1421 => "11111111",
		1422 => "11111111",
		1423 => "11111111",
		1424 => "11111111",
		1425 => "11111111",
		1426 => "11111111",
		1427 => "11111111",
		1428 => "11111111",
		1429 => "11111111",
		1430 => "11111111",
		1431 => "11111111",
		1432 => "11111111",
		1433 => "11111111",
		1434 => "11111111",
		1435 => "11111111",
		1436 => "11111111",
		1437 => "11111111",
		1438 => "11111111",
		1439 => "11111111",
		1440 => "11111111",
		1441 => "11111111",
		1442 => "11111111",
		1443 => "11111111",
		1444 => "11111111",
		1445 => "11111111",
		1446 => "11111111",
		1447 => "11111111",
		1448 => "11111111",
		1449 => "11011100",
		1450 => "01101010",
		1451 => "01101010",
		1452 => "01001101",
		1453 => "11101110",
		1454 => "11111111",
		1455 => "11111111",
		1456 => "11111111",
		1457 => "11111111",
		1458 => "11111111",
		1459 => "11111111",
		1460 => "11111111",
		1461 => "11111001",
		1462 => "01101010",
		1463 => "01100100",
		1464 => "01100100",
		1465 => "01000111",
		1466 => "01111100",
		1467 => "11010111",
		1468 => "11111111",
		1469 => "11101110",
		1470 => "01011001",
		1471 => "11111111",
		1472 => "11111111",
		1473 => "11111111",
		1474 => "11111111",
		1475 => "11111111",
		1476 => "11111111",
		1477 => "11111111",
		1478 => "11111111",
		1479 => "11111111",
		1480 => "11111111",
		1481 => "11111111",
		1482 => "10011110",
		1483 => "01000111",
		1484 => "11000000",
		1485 => "11111111",
		1486 => "11111111",
		1487 => "11111111",
		1488 => "11111111",
		1489 => "11111111",
		1490 => "11111111",
		1491 => "01000111",
		1492 => "01100100",
		1493 => "11111111",
		1494 => "11111111",
		1495 => "11111111",
		1496 => "11111111",
		1497 => "11111111",
		1498 => "11010111",
		1499 => "01001101",
		1500 => "10000001",
		1501 => "11100010",
		1502 => "11111111",
		1503 => "11111111",
		1504 => "11111111",
		1505 => "11111111",
		1506 => "11111111",
		1507 => "11111111",
		1508 => "11111111",
		1509 => "11111111",
		1510 => "11111111",
		1511 => "11111111",
		1512 => "11111111",
		1513 => "11111111",
		1514 => "11111111",
		1515 => "11111111",
		1516 => "11111111",
		1517 => "11111111",
		1518 => "11111111",
		1519 => "11111111",
		1520 => "11111111",
		1521 => "11111111",
		1522 => "11111111",
		1523 => "11111111",
		1524 => "11111111",
		1525 => "11111111",
		1526 => "11111111",
		1527 => "11111111",
		1528 => "11111111",
		1529 => "11111111",
		1530 => "11111111",
		1531 => "11111111",
		1532 => "11111111",
		1533 => "11111111",
		1534 => "11111111",
		1535 => "11111111",
		1536 => "11111111",
		1537 => "11111111",
		1538 => "11111111",
		1539 => "11111111",
		1540 => "11111111",
		1541 => "11111111",
		1542 => "11111111",
		1543 => "11111111",
		1544 => "11111111",
		1545 => "11111111",
		1546 => "11111111",
		1547 => "11111111",
		1548 => "11111111",
		1549 => "11111111",
		1550 => "11111111",
		1551 => "11111111",
		1552 => "11111111",
		1553 => "11111111",
		1554 => "11111111",
		1555 => "11111111",
		1556 => "11111111",
		1557 => "11111111",
		1558 => "11111111",
		1559 => "11111111",
		1560 => "11111111",
		1561 => "11111111",
		1562 => "11111111",
		1563 => "11111111",
		1564 => "11111111",
		1565 => "11111111",
		1566 => "11111111",
		1567 => "11111111",
		1568 => "11111111",
		1569 => "11011100",
		1570 => "10000111",
		1571 => "11011100",
		1572 => "11111111",
		1573 => "11111111",
		1574 => "11111111",
		1575 => "11111111",
		1576 => "11111111",
		1577 => "11101000",
		1578 => "01011110",
		1579 => "11000101",
		1580 => "01000111",
		1581 => "10011000",
		1582 => "11111111",
		1583 => "11111111",
		1584 => "11111111",
		1585 => "11111111",
		1586 => "11111111",
		1587 => "11111111",
		1588 => "11111111",
		1589 => "11000000",
		1590 => "11110011",
		1591 => "11111111",
		1592 => "11101110",
		1593 => "01000111",
		1594 => "01111100",
		1595 => "11111111",
		1596 => "11111111",
		1597 => "11111111",
		1598 => "11000000",
		1599 => "11111111",
		1600 => "11111111",
		1601 => "11111111",
		1602 => "11111111",
		1603 => "11111111",
		1604 => "11111111",
		1605 => "11111111",
		1606 => "11111111",
		1607 => "11111111",
		1608 => "11111111",
		1609 => "11111111",
		1610 => "01101010",
		1611 => "01001101",
		1612 => "11110011",
		1613 => "11111111",
		1614 => "11111111",
		1615 => "11111111",
		1616 => "11111111",
		1617 => "11111111",
		1618 => "11110011",
		1619 => "01000111",
		1620 => "01110101",
		1621 => "11111111",
		1622 => "11111111",
		1623 => "11111111",
		1624 => "11111111",
		1625 => "11111111",
		1626 => "11101000",
		1627 => "01001101",
		1628 => "01010011",
		1629 => "01110101",
		1630 => "11111111",
		1631 => "11111111",
		1632 => "11111111",
		1633 => "11111111",
		1634 => "11111111",
		1635 => "11111111",
		1636 => "11111111",
		1637 => "11111111",
		1638 => "11111111",
		1639 => "11111111",
		1640 => "11111111",
		1641 => "11111111",
		1642 => "11111111",
		1643 => "11111111",
		1644 => "11111111",
		1645 => "11111111",
		1646 => "11111111",
		1647 => "11111111",
		1648 => "11111111",
		1649 => "11111111",
		1650 => "11111111",
		1651 => "11111111",
		1652 => "11111111",
		1653 => "11111111",
		1654 => "11111111",
		1655 => "11111111",
		1656 => "11111111",
		1657 => "11111111",
		1658 => "11111111",
		1659 => "11111111",
		1660 => "11111111",
		1661 => "11111111",
		1662 => "11111111",
		1663 => "11111111",
		1664 => "11111111",
		1665 => "11111111",
		1666 => "11111111",
		1667 => "11111111",
		1668 => "11111111",
		1669 => "11111111",
		1670 => "11111111",
		1671 => "11111111",
		1672 => "11111111",
		1673 => "11111111",
		1674 => "11111111",
		1675 => "11111111",
		1676 => "11111111",
		1677 => "11111111",
		1678 => "11111111",
		1679 => "11111111",
		1680 => "11111111",
		1681 => "11111111",
		1682 => "11111111",
		1683 => "11111111",
		1684 => "11111111",
		1685 => "11111111",
		1686 => "11111111",
		1687 => "11111111",
		1688 => "11111111",
		1689 => "11111111",
		1690 => "11111111",
		1691 => "11111111",
		1692 => "11111111",
		1693 => "11111111",
		1694 => "11111111",
		1695 => "11111111",
		1696 => "11101110",
		1697 => "10011110",
		1698 => "01010011",
		1699 => "01001101",
		1700 => "01001101",
		1701 => "10111010",
		1702 => "11111111",
		1703 => "11111111",
		1704 => "11111111",
		1705 => "11111111",
		1706 => "01000111",
		1707 => "11111111",
		1708 => "11000101",
		1709 => "01000111",
		1710 => "10011000",
		1711 => "11111111",
		1712 => "11111111",
		1713 => "11111111",
		1714 => "11111111",
		1715 => "11111111",
		1716 => "11101110",
		1717 => "01001101",
		1718 => "11111111",
		1719 => "11111111",
		1720 => "11111111",
		1721 => "01110000",
		1722 => "01001101",
		1723 => "11111111",
		1724 => "11111111",
		1725 => "11111111",
		1726 => "11111111",
		1727 => "10011000",
		1728 => "10001100",
		1729 => "11111111",
		1730 => "11111111",
		1731 => "11111111",
		1732 => "11111111",
		1733 => "11111111",
		1734 => "11111111",
		1735 => "11111111",
		1736 => "11111111",
		1737 => "11111111",
		1738 => "01000111",
		1739 => "10101110",
		1740 => "11111111",
		1741 => "11111111",
		1742 => "11111111",
		1743 => "11111111",
		1744 => "11111111",
		1745 => "11111111",
		1746 => "10000001",
		1747 => "01000111",
		1748 => "11000101",
		1749 => "11111111",
		1750 => "11111111",
		1751 => "11111111",
		1752 => "11111111",
		1753 => "11011100",
		1754 => "01000111",
		1755 => "01101010",
		1756 => "11111001",
		1757 => "11111111",
		1758 => "11111111",
		1759 => "11111111",
		1760 => "11111111",
		1761 => "11111111",
		1762 => "11111111",
		1763 => "11111111",
		1764 => "11111111",
		1765 => "11111111",
		1766 => "11111111",
		1767 => "11111111",
		1768 => "11111111",
		1769 => "11111111",
		1770 => "11111111",
		1771 => "11111111",
		1772 => "11111111",
		1773 => "11111111",
		1774 => "11111111",
		1775 => "11111111",
		1776 => "11111111",
		1777 => "11111111",
		1778 => "11111111",
		1779 => "11111111",
		1780 => "11111111",
		1781 => "11111111",
		1782 => "11111111",
		1783 => "11111111",
		1784 => "11111111",
		1785 => "11111111",
		1786 => "11111111",
		1787 => "11111111",
		1788 => "11111111",
		1789 => "11111111",
		1790 => "11111111",
		1791 => "11111111",
		1792 => "11111111",
		1793 => "11111111",
		1794 => "11111111",
		1795 => "11111111",
		1796 => "11111111",
		1797 => "11111111",
		1798 => "11111111",
		1799 => "11111111",
		1800 => "11111111",
		1801 => "11111111",
		1802 => "11111111",
		1803 => "11111111",
		1804 => "11111111",
		1805 => "11111111",
		1806 => "11111111",
		1807 => "11111111",
		1808 => "11111111",
		1809 => "11111111",
		1810 => "11111111",
		1811 => "11111111",
		1812 => "11111111",
		1813 => "11111111",
		1814 => "11111111",
		1815 => "11111111",
		1816 => "11111111",
		1817 => "11111111",
		1818 => "11111111",
		1819 => "11111111",
		1820 => "11111111",
		1821 => "11111111",
		1822 => "11111111",
		1823 => "11111111",
		1824 => "11111111",
		1825 => "11111001",
		1826 => "01011001",
		1827 => "10101110",
		1828 => "01010011",
		1829 => "01000111",
		1830 => "10101001",
		1831 => "11111111",
		1832 => "11111111",
		1833 => "11111111",
		1834 => "01011001",
		1835 => "11101000",
		1836 => "11111111",
		1837 => "01101010",
		1838 => "01001101",
		1839 => "11101110",
		1840 => "11111111",
		1841 => "11111111",
		1842 => "11111111",
		1843 => "11111111",
		1844 => "10101001",
		1845 => "10000111",
		1846 => "11111111",
		1847 => "11111111",
		1848 => "11111111",
		1849 => "10000111",
		1850 => "01000111",
		1851 => "11101110",
		1852 => "11111111",
		1853 => "11010111",
		1854 => "11010001",
		1855 => "01011001",
		1856 => "10001100",
		1857 => "11111111",
		1858 => "11111111",
		1859 => "11111111",
		1860 => "11111111",
		1861 => "11111111",
		1862 => "11111111",
		1863 => "11111111",
		1864 => "11111111",
		1865 => "11111111",
		1866 => "01000111",
		1867 => "11100010",
		1868 => "11111111",
		1869 => "11111111",
		1870 => "11111111",
		1871 => "11111111",
		1872 => "11111111",
		1873 => "11011100",
		1874 => "01000111",
		1875 => "01101010",
		1876 => "11111111",
		1877 => "11111111",
		1878 => "11111111",
		1879 => "11111111",
		1880 => "11111111",
		1881 => "10000001",
		1882 => "01000111",
		1883 => "11000101",
		1884 => "11111111",
		1885 => "11111111",
		1886 => "11111111",
		1887 => "11111111",
		1888 => "11111111",
		1889 => "11111111",
		1890 => "11111111",
		1891 => "11111111",
		1892 => "11111111",
		1893 => "11111111",
		1894 => "11111111",
		1895 => "11111111",
		1896 => "11111111",
		1897 => "11111111",
		1898 => "11111111",
		1899 => "11111111",
		1900 => "11111111",
		1901 => "11111111",
		1902 => "11111111",
		1903 => "11111111",
		1904 => "11111111",
		1905 => "11111111",
		1906 => "11111111",
		1907 => "11111111",
		1908 => "11111111",
		1909 => "11111111",
		1910 => "11111111",
		1911 => "11111111",
		1912 => "11111111",
		1913 => "11111111",
		1914 => "11111111",
		1915 => "11111111",
		1916 => "11111111",
		1917 => "11111111",
		1918 => "11111111",
		1919 => "11111111",
		1920 => "11111111",
		1921 => "11111111",
		1922 => "11111111",
		1923 => "11111111",
		1924 => "11111111",
		1925 => "11111111",
		1926 => "11111111",
		1927 => "11111111",
		1928 => "11111111",
		1929 => "11111111",
		1930 => "11111111",
		1931 => "11111111",
		1932 => "11111111",
		1933 => "11111111",
		1934 => "11111111",
		1935 => "11111111",
		1936 => "11111111",
		1937 => "11111111",
		1938 => "11111111",
		1939 => "11111111",
		1940 => "11111111",
		1941 => "11111111",
		1942 => "11111111",
		1943 => "11111111",
		1944 => "11111111",
		1945 => "11111111",
		1946 => "11111111",
		1947 => "11111111",
		1948 => "11111111",
		1949 => "11111111",
		1950 => "11111111",
		1951 => "11111111",
		1952 => "11111111",
		1953 => "11111111",
		1954 => "10101110",
		1955 => "10000001",
		1956 => "11011100",
		1957 => "01011110",
		1958 => "01000111",
		1959 => "10010011",
		1960 => "11111111",
		1961 => "11111111",
		1962 => "01011110",
		1963 => "11100010",
		1964 => "11111111",
		1965 => "11000101",
		1966 => "01000111",
		1967 => "10011000",
		1968 => "11111111",
		1969 => "11111111",
		1970 => "11111111",
		1971 => "11111111",
		1972 => "01100100",
		1973 => "10101110",
		1974 => "11111111",
		1975 => "11111111",
		1976 => "11000000",
		1977 => "01011001",
		1978 => "01000111",
		1979 => "01001101",
		1980 => "01110101",
		1981 => "10000001",
		1982 => "10100011",
		1983 => "10110100",
		1984 => "11100010",
		1985 => "11111111",
		1986 => "11111111",
		1987 => "11111111",
		1988 => "11111111",
		1989 => "11111111",
		1990 => "11111111",
		1991 => "11111111",
		1992 => "10111010",
		1993 => "10001100",
		1994 => "01011110",
		1995 => "11111111",
		1996 => "11111111",
		1997 => "11111111",
		1998 => "11111111",
		1999 => "11111111",
		2000 => "11011100",
		2001 => "01011110",
		2002 => "01000111",
		2003 => "11001011",
		2004 => "11111111",
		2005 => "11111111",
		2006 => "11111111",
		2007 => "11111111",
		2008 => "11010001",
		2009 => "01000111",
		2010 => "01101010",
		2011 => "11111111",
		2012 => "11111111",
		2013 => "11111111",
		2014 => "11111111",
		2015 => "11111111",
		2016 => "11111111",
		2017 => "11111111",
		2018 => "11111111",
		2019 => "11111111",
		2020 => "11111111",
		2021 => "11111111",
		2022 => "11111111",
		2023 => "11111111",
		2024 => "11111111",
		2025 => "11111111",
		2026 => "11111111",
		2027 => "11111111",
		2028 => "11111111",
		2029 => "11111111",
		2030 => "11111111",
		2031 => "11111111",
		2032 => "11111111",
		2033 => "11111111",
		2034 => "11111111",
		2035 => "11111111",
		2036 => "11111111",
		2037 => "11111111",
		2038 => "11111111",
		2039 => "11111111",
		2040 => "11111111",
		2041 => "11111111",
		2042 => "11111111",
		2043 => "11111111",
		2044 => "11111111",
		2045 => "11111111",
		2046 => "11111111",
		2047 => "11111111",
		2048 => "11111111",
		2049 => "11111111",
		2050 => "11111111",
		2051 => "11111111",
		2052 => "11111111",
		2053 => "11111111",
		2054 => "11111111",
		2055 => "11111111",
		2056 => "11111111",
		2057 => "11111111",
		2058 => "11111111",
		2059 => "11111111",
		2060 => "11111111",
		2061 => "11111111",
		2062 => "11111111",
		2063 => "11111111",
		2064 => "11111111",
		2065 => "11111111",
		2066 => "11111111",
		2067 => "11111111",
		2068 => "11111111",
		2069 => "11111111",
		2070 => "11111111",
		2071 => "11111111",
		2072 => "11111111",
		2073 => "11111111",
		2074 => "11111111",
		2075 => "11000000",
		2076 => "10011110",
		2077 => "11111111",
		2078 => "11111111",
		2079 => "11111111",
		2080 => "11111111",
		2081 => "11111111",
		2082 => "11111001",
		2083 => "01011001",
		2084 => "11011100",
		2085 => "11101000",
		2086 => "01101010",
		2087 => "01000111",
		2088 => "10000111",
		2089 => "11111001",
		2090 => "01110101",
		2091 => "11010001",
		2092 => "11111111",
		2093 => "11111111",
		2094 => "01101010",
		2095 => "01001101",
		2096 => "11101110",
		2097 => "11111111",
		2098 => "11101000",
		2099 => "01110101",
		2100 => "01000111",
		2101 => "01011110",
		2102 => "11111111",
		2103 => "11111111",
		2104 => "11010111",
		2105 => "11010001",
		2106 => "11111111",
		2107 => "11111111",
		2108 => "11111111",
		2109 => "11111111",
		2110 => "11111111",
		2111 => "11111111",
		2112 => "11111111",
		2113 => "11111111",
		2114 => "11111111",
		2115 => "11111111",
		2116 => "11111111",
		2117 => "11111111",
		2118 => "11111111",
		2119 => "11111111",
		2120 => "11111001",
		2121 => "11000101",
		2122 => "01101010",
		2123 => "01111100",
		2124 => "10100011",
		2125 => "11000000",
		2126 => "11001011",
		2127 => "10011000",
		2128 => "01010011",
		2129 => "01100100",
		2130 => "11010111",
		2131 => "11111111",
		2132 => "11111111",
		2133 => "11111111",
		2134 => "11111111",
		2135 => "11111111",
		2136 => "01101010",
		2137 => "01000111",
		2138 => "11010111",
		2139 => "11111111",
		2140 => "11111111",
		2141 => "11111111",
		2142 => "11111111",
		2143 => "11101000",
		2144 => "10101001",
		2145 => "01110000",
		2146 => "01000111",
		2147 => "01101010",
		2148 => "10000001",
		2149 => "11010111",
		2150 => "11111111",
		2151 => "11111111",
		2152 => "11111111",
		2153 => "11111111",
		2154 => "11111111",
		2155 => "11111111",
		2156 => "11111111",
		2157 => "11111111",
		2158 => "11111111",
		2159 => "11111111",
		2160 => "11111111",
		2161 => "11111111",
		2162 => "11111111",
		2163 => "11111111",
		2164 => "11111111",
		2165 => "11111111",
		2166 => "11111111",
		2167 => "11111111",
		2168 => "11111111",
		2169 => "11111111",
		2170 => "11111111",
		2171 => "11111111",
		2172 => "11111111",
		2173 => "11111111",
		2174 => "11111111",
		2175 => "11111111",
		2176 => "11111111",
		2177 => "11111111",
		2178 => "11111111",
		2179 => "11111111",
		2180 => "11111111",
		2181 => "11111111",
		2182 => "11111111",
		2183 => "11111111",
		2184 => "11111111",
		2185 => "11111111",
		2186 => "11111111",
		2187 => "11111111",
		2188 => "11111111",
		2189 => "11111111",
		2190 => "11111111",
		2191 => "11111111",
		2192 => "11111111",
		2193 => "11111111",
		2194 => "11111111",
		2195 => "11111111",
		2196 => "11111111",
		2197 => "11111111",
		2198 => "11111111",
		2199 => "11111111",
		2200 => "11111111",
		2201 => "11111111",
		2202 => "10101001",
		2203 => "01101010",
		2204 => "01001101",
		2205 => "10101001",
		2206 => "11111111",
		2207 => "11111111",
		2208 => "11111111",
		2209 => "11111111",
		2210 => "11111111",
		2211 => "10101110",
		2212 => "10000001",
		2213 => "11111111",
		2214 => "11110011",
		2215 => "01110101",
		2216 => "01000111",
		2217 => "01110101",
		2218 => "01101010",
		2219 => "11000101",
		2220 => "11111111",
		2221 => "11111111",
		2222 => "11000101",
		2223 => "01000111",
		2224 => "01100100",
		2225 => "01100100",
		2226 => "11010011",
		2227 => "11100010",
		2228 => "11111111",
		2229 => "11111111",
		2230 => "11111111",
		2231 => "11111111",
		2232 => "11111111",
		2233 => "11111111",
		2234 => "11111111",
		2235 => "11111111",
		2236 => "11111111",
		2237 => "11111111",
		2238 => "11111111",
		2239 => "11111111",
		2240 => "11111111",
		2241 => "11111111",
		2242 => "11111111",
		2243 => "11111111",
		2244 => "11111111",
		2245 => "11111111",
		2246 => "11111111",
		2247 => "11111111",
		2248 => "11111111",
		2249 => "11111111",
		2250 => "11111111",
		2251 => "11101000",
		2252 => "10110100",
		2253 => "10100011",
		2254 => "01110101",
		2255 => "10001100",
		2256 => "10101110",
		2257 => "11111001",
		2258 => "11111111",
		2259 => "11111111",
		2260 => "11111111",
		2261 => "11111111",
		2262 => "11111111",
		2263 => "11000101",
		2264 => "01000111",
		2265 => "10000001",
		2266 => "11111111",
		2267 => "11111111",
		2268 => "11111111",
		2269 => "11111111",
		2270 => "11001011",
		2271 => "01010011",
		2272 => "01000111",
		2273 => "01101010",
		2274 => "10101110",
		2275 => "11000000",
		2276 => "10100011",
		2277 => "01101010",
		2278 => "10010011",
		2279 => "11110011",
		2280 => "11111111",
		2281 => "11111111",
		2282 => "11111111",
		2283 => "11111111",
		2284 => "11111111",
		2285 => "11111111",
		2286 => "11111111",
		2287 => "11111111",
		2288 => "11111111",
		2289 => "11111111",
		2290 => "11111111",
		2291 => "11111111",
		2292 => "11111111",
		2293 => "11111111",
		2294 => "11111111",
		2295 => "11111111",
		2296 => "11111111",
		2297 => "11111111",
		2298 => "11111111",
		2299 => "11111111",
		2300 => "11111111",
		2301 => "11111111",
		2302 => "11111111",
		2303 => "11111111",
		2304 => "11111111",
		2305 => "11111111",
		2306 => "11111111",
		2307 => "11111111",
		2308 => "11111111",
		2309 => "11111111",
		2310 => "11111111",
		2311 => "11111111",
		2312 => "11111111",
		2313 => "11111111",
		2314 => "11111111",
		2315 => "11111111",
		2316 => "11111111",
		2317 => "11111111",
		2318 => "11111111",
		2319 => "11111111",
		2320 => "11111111",
		2321 => "11111111",
		2322 => "11111111",
		2323 => "11111111",
		2324 => "11111111",
		2325 => "11111111",
		2326 => "11111111",
		2327 => "11111111",
		2328 => "11111111",
		2329 => "10010011",
		2330 => "10011110",
		2331 => "11111111",
		2332 => "11101110",
		2333 => "10110100",
		2334 => "11111111",
		2335 => "11111111",
		2336 => "11111111",
		2337 => "11111111",
		2338 => "11111111",
		2339 => "11111001",
		2340 => "01011001",
		2341 => "11011100",
		2342 => "11111111",
		2343 => "11111001",
		2344 => "10000111",
		2345 => "01000111",
		2346 => "01000111",
		2347 => "10111010",
		2348 => "11111111",
		2349 => "11111111",
		2350 => "10001100",
		2351 => "01011110",
		2352 => "10110100",
		2353 => "11111001",
		2354 => "11111111",
		2355 => "11111111",
		2356 => "11111111",
		2357 => "11111111",
		2358 => "11111111",
		2359 => "11111111",
		2360 => "11111111",
		2361 => "11111111",
		2362 => "11111111",
		2363 => "11111111",
		2364 => "11111111",
		2365 => "11111111",
		2366 => "11111111",
		2367 => "11111111",
		2368 => "11111111",
		2369 => "11111111",
		2370 => "11111111",
		2371 => "11111111",
		2372 => "11111111",
		2373 => "11111111",
		2374 => "11111111",
		2375 => "11111111",
		2376 => "11111111",
		2377 => "11111111",
		2378 => "11111111",
		2379 => "11111111",
		2380 => "11111111",
		2381 => "11111111",
		2382 => "11111111",
		2383 => "11111111",
		2384 => "11111111",
		2385 => "11111111",
		2386 => "11111111",
		2387 => "11111111",
		2388 => "11111111",
		2389 => "11111111",
		2390 => "11111111",
		2391 => "01101010",
		2392 => "01000111",
		2393 => "11011100",
		2394 => "11111111",
		2395 => "11111111",
		2396 => "11111111",
		2397 => "11111111",
		2398 => "01000111",
		2399 => "01001101",
		2400 => "11000000",
		2401 => "11111111",
		2402 => "11111111",
		2403 => "11111111",
		2404 => "11111111",
		2405 => "11111111",
		2406 => "10101110",
		2407 => "01110000",
		2408 => "11101000",
		2409 => "11111111",
		2410 => "11111111",
		2411 => "11111111",
		2412 => "11111111",
		2413 => "11111111",
		2414 => "11111111",
		2415 => "11111111",
		2416 => "11111111",
		2417 => "11111111",
		2418 => "11111111",
		2419 => "11111111",
		2420 => "11111111",
		2421 => "11111111",
		2422 => "11111111",
		2423 => "11111111",
		2424 => "11111111",
		2425 => "11111111",
		2426 => "11111111",
		2427 => "11111111",
		2428 => "11111111",
		2429 => "11111111",
		2430 => "11111111",
		2431 => "11111111",
		2432 => "11111111",
		2433 => "11111111",
		2434 => "11111111",
		2435 => "11111111",
		2436 => "11111111",
		2437 => "11111111",
		2438 => "11111111",
		2439 => "11111111",
		2440 => "11111111",
		2441 => "11111111",
		2442 => "11111111",
		2443 => "11111111",
		2444 => "11111111",
		2445 => "11111111",
		2446 => "11111111",
		2447 => "11111111",
		2448 => "11111111",
		2449 => "11111111",
		2450 => "11111111",
		2451 => "11111111",
		2452 => "11111111",
		2453 => "11111111",
		2454 => "11111111",
		2455 => "11110011",
		2456 => "10000001",
		2457 => "10111010",
		2458 => "11111111",
		2459 => "11111111",
		2460 => "11111111",
		2461 => "11111111",
		2462 => "11110011",
		2463 => "11111111",
		2464 => "11111111",
		2465 => "11111111",
		2466 => "11111111",
		2467 => "11111111",
		2468 => "10101110",
		2469 => "10000001",
		2470 => "11111111",
		2471 => "11111111",
		2472 => "11111111",
		2473 => "10011000",
		2474 => "01000111",
		2475 => "10101001",
		2476 => "11111111",
		2477 => "11101000",
		2478 => "10111010",
		2479 => "11111111",
		2480 => "11111111",
		2481 => "11111111",
		2482 => "11111111",
		2483 => "11111111",
		2484 => "11111111",
		2485 => "11111111",
		2486 => "11111111",
		2487 => "11111111",
		2488 => "11111111",
		2489 => "11111111",
		2490 => "11111111",
		2491 => "11111111",
		2492 => "11111111",
		2493 => "11111111",
		2494 => "11111111",
		2495 => "11111111",
		2496 => "11111111",
		2497 => "11111111",
		2498 => "11111111",
		2499 => "11111111",
		2500 => "11111111",
		2501 => "11111111",
		2502 => "11111111",
		2503 => "11111111",
		2504 => "11111111",
		2505 => "11111111",
		2506 => "11111111",
		2507 => "11111111",
		2508 => "11111111",
		2509 => "11111111",
		2510 => "11111111",
		2511 => "11111111",
		2512 => "11111111",
		2513 => "11111111",
		2514 => "11111111",
		2515 => "11111111",
		2516 => "11101110",
		2517 => "11011100",
		2518 => "10101110",
		2519 => "01000111",
		2520 => "10010011",
		2521 => "11111111",
		2522 => "11111111",
		2523 => "11111111",
		2524 => "11111111",
		2525 => "11101110",
		2526 => "01001101",
		2527 => "11001011",
		2528 => "11111111",
		2529 => "11111111",
		2530 => "11111111",
		2531 => "11111111",
		2532 => "11111111",
		2533 => "11111111",
		2534 => "11111111",
		2535 => "11001011",
		2536 => "01101010",
		2537 => "11110011",
		2538 => "11111111",
		2539 => "11111111",
		2540 => "11111111",
		2541 => "11111111",
		2542 => "11111111",
		2543 => "11111111",
		2544 => "11111111",
		2545 => "11111111",
		2546 => "11111111",
		2547 => "11111111",
		2548 => "11111111",
		2549 => "11111111",
		2550 => "11111111",
		2551 => "11111111",
		2552 => "11111111",
		2553 => "11111111",
		2554 => "11111111",
		2555 => "11111111",
		2556 => "11111111",
		2557 => "11111111",
		2558 => "11111111",
		2559 => "11111111",
		2560 => "11111111",
		2561 => "11111111",
		2562 => "11111111",
		2563 => "11111111",
		2564 => "11111111",
		2565 => "11111111",
		2566 => "11111111",
		2567 => "11111111",
		2568 => "11111111",
		2569 => "11111111",
		2570 => "11111111",
		2571 => "11111111",
		2572 => "11111111",
		2573 => "11111111",
		2574 => "11111111",
		2575 => "11111111",
		2576 => "11111111",
		2577 => "11111111",
		2578 => "11111111",
		2579 => "11111111",
		2580 => "11111111",
		2581 => "11111111",
		2582 => "11101110",
		2583 => "01101010",
		2584 => "01110000",
		2585 => "11111111",
		2586 => "11111111",
		2587 => "11111111",
		2588 => "11111111",
		2589 => "11101110",
		2590 => "01110000",
		2591 => "11110011",
		2592 => "11111111",
		2593 => "11111111",
		2594 => "11111111",
		2595 => "11111111",
		2596 => "11111001",
		2597 => "01011001",
		2598 => "11011100",
		2599 => "11111111",
		2600 => "11111111",
		2601 => "11111111",
		2602 => "10101110",
		2603 => "10100011",
		2604 => "11111111",
		2605 => "11111111",
		2606 => "11111111",
		2607 => "11111111",
		2608 => "11111111",
		2609 => "11111111",
		2610 => "11111111",
		2611 => "11111111",
		2612 => "11111111",
		2613 => "11111111",
		2614 => "11111111",
		2615 => "11111111",
		2616 => "11111111",
		2617 => "11111111",
		2618 => "11111111",
		2619 => "11111111",
		2620 => "11111111",
		2621 => "11111111",
		2622 => "11111111",
		2623 => "11111111",
		2624 => "11111111",
		2625 => "11111111",
		2626 => "11111111",
		2627 => "11111111",
		2628 => "11111111",
		2629 => "11111111",
		2630 => "11111111",
		2631 => "11111111",
		2632 => "11111111",
		2633 => "11111111",
		2634 => "11111111",
		2635 => "11111111",
		2636 => "11111111",
		2637 => "11111111",
		2638 => "11111111",
		2639 => "11111111",
		2640 => "11111111",
		2641 => "11111111",
		2642 => "11111111",
		2643 => "11111111",
		2644 => "11011100",
		2645 => "01110101",
		2646 => "01000111",
		2647 => "01000111",
		2648 => "11101110",
		2649 => "11111111",
		2650 => "11111111",
		2651 => "11111111",
		2652 => "11111111",
		2653 => "10000111",
		2654 => "10100011",
		2655 => "11111111",
		2656 => "11111111",
		2657 => "11111111",
		2658 => "11111111",
		2659 => "11111111",
		2660 => "11111111",
		2661 => "11111111",
		2662 => "11111111",
		2663 => "11101000",
		2664 => "01000111",
		2665 => "10101001",
		2666 => "11111111",
		2667 => "11111111",
		2668 => "11111111",
		2669 => "11111111",
		2670 => "11111111",
		2671 => "11111111",
		2672 => "11111111",
		2673 => "11111111",
		2674 => "11111111",
		2675 => "11111111",
		2676 => "11111111",
		2677 => "11111111",
		2678 => "11111111",
		2679 => "11111111",
		2680 => "11111111",
		2681 => "11111111",
		2682 => "11111111",
		2683 => "11111111",
		2684 => "11111111",
		2685 => "11111111",
		2686 => "11111111",
		2687 => "11111111",
		2688 => "11111111",
		2689 => "11111111",
		2690 => "11111111",
		2691 => "11111111",
		2692 => "11111111",
		2693 => "11111111",
		2694 => "11111111",
		2695 => "11111111",
		2696 => "11111111",
		2697 => "11111111",
		2698 => "11111111",
		2699 => "11111111",
		2700 => "11111111",
		2701 => "11111111",
		2702 => "11111111",
		2703 => "11111111",
		2704 => "11111111",
		2705 => "11111111",
		2706 => "11111111",
		2707 => "11111111",
		2708 => "11111111",
		2709 => "11011100",
		2710 => "01011110",
		2711 => "01011110",
		2712 => "01000111",
		2713 => "10001100",
		2714 => "11111111",
		2715 => "11111111",
		2716 => "11111111",
		2717 => "11111111",
		2718 => "01111100",
		2719 => "01110101",
		2720 => "11111001",
		2721 => "11111111",
		2722 => "11111111",
		2723 => "11111111",
		2724 => "11111111",
		2725 => "10101110",
		2726 => "01111100",
		2727 => "11010001",
		2728 => "11100010",
		2729 => "11111111",
		2730 => "11111111",
		2731 => "11111111",
		2732 => "11111111",
		2733 => "11111111",
		2734 => "11111111",
		2735 => "11111111",
		2736 => "11111111",
		2737 => "11111111",
		2738 => "11111111",
		2739 => "11111111",
		2740 => "11111111",
		2741 => "11111111",
		2742 => "11111111",
		2743 => "11111111",
		2744 => "11111111",
		2745 => "11111111",
		2746 => "11111111",
		2747 => "11111111",
		2748 => "11111111",
		2749 => "11111111",
		2750 => "11111111",
		2751 => "11111111",
		2752 => "11111111",
		2753 => "11111111",
		2754 => "11111111",
		2755 => "11111111",
		2756 => "11111111",
		2757 => "11111111",
		2758 => "11111111",
		2759 => "11111111",
		2760 => "11111111",
		2761 => "11111111",
		2762 => "11111111",
		2763 => "11111111",
		2764 => "11111111",
		2765 => "11111111",
		2766 => "11111111",
		2767 => "11111111",
		2768 => "11111111",
		2769 => "11111111",
		2770 => "11111111",
		2771 => "11111111",
		2772 => "11111111",
		2773 => "11111111",
		2774 => "11010001",
		2775 => "01110000",
		2776 => "10011000",
		2777 => "11111111",
		2778 => "11111111",
		2779 => "11111111",
		2780 => "11111111",
		2781 => "01010011",
		2782 => "11111001",
		2783 => "11111111",
		2784 => "11111111",
		2785 => "11111111",
		2786 => "11111111",
		2787 => "11111111",
		2788 => "11111111",
		2789 => "11111111",
		2790 => "11111111",
		2791 => "10101001",
		2792 => "01110101",
		2793 => "11111001",
		2794 => "11111111",
		2795 => "11111111",
		2796 => "11111111",
		2797 => "11111111",
		2798 => "11111111",
		2799 => "11111111",
		2800 => "11111111",
		2801 => "11111111",
		2802 => "11111111",
		2803 => "11111111",
		2804 => "11111111",
		2805 => "11111111",
		2806 => "11111111",
		2807 => "11111111",
		2808 => "11111111",
		2809 => "11111111",
		2810 => "11111111",
		2811 => "11111111",
		2812 => "11111111",
		2813 => "11111111",
		2814 => "11111111",
		2815 => "11111111",
		2816 => "11111111",
		2817 => "11111111",
		2818 => "11111111",
		2819 => "11111111",
		2820 => "11111111",
		2821 => "11111111",
		2822 => "11111111",
		2823 => "11111111",
		2824 => "11111111",
		2825 => "11111111",
		2826 => "11111111",
		2827 => "11111111",
		2828 => "11111111",
		2829 => "11111111",
		2830 => "11111111",
		2831 => "11111111",
		2832 => "11111111",
		2833 => "11111111",
		2834 => "11111111",
		2835 => "11111111",
		2836 => "11111111",
		2837 => "11101110",
		2838 => "11111001",
		2839 => "11110011",
		2840 => "01011110",
		2841 => "01000111",
		2842 => "10100011",
		2843 => "11111111",
		2844 => "11111111",
		2845 => "10111010",
		2846 => "01111100",
		2847 => "10000001",
		2848 => "10000001",
		2849 => "11111111",
		2850 => "11111111",
		2851 => "11111111",
		2852 => "11111111",
		2853 => "11000101",
		2854 => "01000111",
		2855 => "10000001",
		2856 => "11011100",
		2857 => "11111111",
		2858 => "11111111",
		2859 => "11111111",
		2860 => "11111111",
		2861 => "11111111",
		2862 => "11111111",
		2863 => "11111111",
		2864 => "11111111",
		2865 => "11111111",
		2866 => "11111111",
		2867 => "11111111",
		2868 => "11111111",
		2869 => "11111111",
		2870 => "11010001",
		2871 => "11010001",
		2872 => "11010001",
		2873 => "11010001",
		2874 => "11010001",
		2875 => "11110011",
		2876 => "11111111",
		2877 => "11111111",
		2878 => "11111111",
		2879 => "11111111",
		2880 => "11111111",
		2881 => "11111111",
		2882 => "11100010",
		2883 => "11010001",
		2884 => "11010001",
		2885 => "11010001",
		2886 => "10101110",
		2887 => "10100011",
		2888 => "10100011",
		2889 => "11000000",
		2890 => "11010001",
		2891 => "11100010",
		2892 => "11111111",
		2893 => "11111111",
		2894 => "11111111",
		2895 => "11111111",
		2896 => "11111111",
		2897 => "11111111",
		2898 => "11111111",
		2899 => "11111111",
		2900 => "11111111",
		2901 => "11111111",
		2902 => "11111111",
		2903 => "11111111",
		2904 => "11001011",
		2905 => "11111111",
		2906 => "11111111",
		2907 => "11111111",
		2908 => "11101110",
		2909 => "01000111",
		2910 => "11111111",
		2911 => "11111111",
		2912 => "11111111",
		2913 => "11111111",
		2914 => "11111111",
		2915 => "11111111",
		2916 => "11111111",
		2917 => "11111111",
		2918 => "11111111",
		2919 => "11001011",
		2920 => "11110011",
		2921 => "11111111",
		2922 => "11111111",
		2923 => "11111111",
		2924 => "11111111",
		2925 => "11111111",
		2926 => "11111111",
		2927 => "11111111",
		2928 => "11111111",
		2929 => "11111111",
		2930 => "11111111",
		2931 => "11111111",
		2932 => "11111111",
		2933 => "11111111",
		2934 => "11111111",
		2935 => "11111111",
		2936 => "11111111",
		2937 => "11111111",
		2938 => "11111111",
		2939 => "11111111",
		2940 => "11111111",
		2941 => "11111111",
		2942 => "11111111",
		2943 => "11111111",
		2944 => "11111111",
		2945 => "11111111",
		2946 => "11111111",
		2947 => "11111111",
		2948 => "11111111",
		2949 => "11111111",
		2950 => "11111111",
		2951 => "11111111",
		2952 => "11111111",
		2953 => "11111111",
		2954 => "11111111",
		2955 => "11111111",
		2956 => "11111111",
		2957 => "11111111",
		2958 => "11111111",
		2959 => "11111111",
		2960 => "11111111",
		2961 => "11111111",
		2962 => "11111111",
		2963 => "11111111",
		2964 => "11111111",
		2965 => "11111111",
		2966 => "11111111",
		2967 => "11111111",
		2968 => "11101000",
		2969 => "01011001",
		2970 => "01000111",
		2971 => "10110100",
		2972 => "10011110",
		2973 => "10010011",
		2974 => "11111111",
		2975 => "11111111",
		2976 => "11110011",
		2977 => "10101001",
		2978 => "11010001",
		2979 => "11111111",
		2980 => "11110011",
		2981 => "10000111",
		2982 => "11011100",
		2983 => "11111111",
		2984 => "11111111",
		2985 => "11111111",
		2986 => "11111111",
		2987 => "11111111",
		2988 => "11111111",
		2989 => "11111111",
		2990 => "11111111",
		2991 => "11111111",
		2992 => "11111111",
		2993 => "11010111",
		2994 => "10101001",
		2995 => "01111100",
		2996 => "01011110",
		2997 => "01000111",
		2998 => "01000111",
		2999 => "01000111",
		3000 => "01000111",
		3001 => "01000111",
		3002 => "01000111",
		3003 => "01000111",
		3004 => "01000111",
		3005 => "01010011",
		3006 => "01110101",
		3007 => "01110101",
		3008 => "01001101",
		3009 => "01000111",
		3010 => "01000111",
		3011 => "01000111",
		3012 => "01000111",
		3013 => "01000111",
		3014 => "01000111",
		3015 => "01000111",
		3016 => "01000111",
		3017 => "01000111",
		3018 => "01000111",
		3019 => "01000111",
		3020 => "01010011",
		3021 => "10000001",
		3022 => "10101001",
		3023 => "11011100",
		3024 => "11111111",
		3025 => "11111111",
		3026 => "11111111",
		3027 => "11111111",
		3028 => "11111111",
		3029 => "11111111",
		3030 => "11111111",
		3031 => "11111111",
		3032 => "11111111",
		3033 => "11111111",
		3034 => "11111111",
		3035 => "11111111",
		3036 => "11110011",
		3037 => "01000111",
		3038 => "11111111",
		3039 => "11111111",
		3040 => "11111111",
		3041 => "11111111",
		3042 => "11101000",
		3043 => "11111111",
		3044 => "11111111",
		3045 => "11111111",
		3046 => "11111111",
		3047 => "11111111",
		3048 => "11111111",
		3049 => "11111111",
		3050 => "11111111",
		3051 => "11111111",
		3052 => "11111111",
		3053 => "11111111",
		3054 => "11111111",
		3055 => "11111111",
		3056 => "11111111",
		3057 => "11111111",
		3058 => "11111111",
		3059 => "11111111",
		3060 => "11111111",
		3061 => "11111111",
		3062 => "11111111",
		3063 => "11111111",
		3064 => "11111111",
		3065 => "11111111",
		3066 => "11111111",
		3067 => "11111111",
		3068 => "11111111",
		3069 => "11111111",
		3070 => "11111111",
		3071 => "11111111",
		3072 => "11111111",
		3073 => "11111111",
		3074 => "11111111",
		3075 => "11111111",
		3076 => "11111111",
		3077 => "11111111",
		3078 => "11111111",
		3079 => "11111111",
		3080 => "11111111",
		3081 => "11111111",
		3082 => "11111111",
		3083 => "11111111",
		3084 => "11111111",
		3085 => "11111111",
		3086 => "11111111",
		3087 => "11111111",
		3088 => "11111111",
		3089 => "11111111",
		3090 => "11111111",
		3091 => "11111111",
		3092 => "11111111",
		3093 => "11111111",
		3094 => "11111111",
		3095 => "11111111",
		3096 => "11111111",
		3097 => "11011100",
		3098 => "01010011",
		3099 => "01000111",
		3100 => "10001100",
		3101 => "11111111",
		3102 => "11111111",
		3103 => "11111111",
		3104 => "11111111",
		3105 => "11000101",
		3106 => "01011001",
		3107 => "11101110",
		3108 => "11111111",
		3109 => "11111111",
		3110 => "11111111",
		3111 => "11111111",
		3112 => "11111111",
		3113 => "11111111",
		3114 => "11111111",
		3115 => "11111111",
		3116 => "11111111",
		3117 => "11111111",
		3118 => "11111111",
		3119 => "10101001",
		3120 => "01010011",
		3121 => "01000111",
		3122 => "01000111",
		3123 => "01100100",
		3124 => "10000001",
		3125 => "10100011",
		3126 => "10100011",
		3127 => "10100011",
		3128 => "10000111",
		3129 => "01011110",
		3130 => "01000111",
		3131 => "01000111",
		3132 => "01000111",
		3133 => "01000111",
		3134 => "01100100",
		3135 => "01110101",
		3136 => "10100011",
		3137 => "10100011",
		3138 => "11000101",
		3139 => "11010001",
		3140 => "11101000",
		3141 => "11111111",
		3142 => "11111111",
		3143 => "11111111",
		3144 => "11111111",
		3145 => "11110011",
		3146 => "11010001",
		3147 => "10111010",
		3148 => "10011110",
		3149 => "01101010",
		3150 => "01000111",
		3151 => "01000111",
		3152 => "10000111",
		3153 => "11111111",
		3154 => "11111111",
		3155 => "11111111",
		3156 => "11111111",
		3157 => "11111111",
		3158 => "11111111",
		3159 => "11111111",
		3160 => "11111111",
		3161 => "11111111",
		3162 => "11111111",
		3163 => "11111111",
		3164 => "11111111",
		3165 => "01110000",
		3166 => "11111111",
		3167 => "11111111",
		3168 => "11111111",
		3169 => "11111111",
		3170 => "10000001",
		3171 => "10101110",
		3172 => "11111111",
		3173 => "11111111",
		3174 => "11111111",
		3175 => "11111111",
		3176 => "11111111",
		3177 => "11111111",
		3178 => "11111111",
		3179 => "11111111",
		3180 => "11111111",
		3181 => "11010111",
		3182 => "11010001",
		3183 => "11111111",
		3184 => "11111111",
		3185 => "11111111",
		3186 => "11111111",
		3187 => "11111111",
		3188 => "11111111",
		3189 => "11111111",
		3190 => "11111111",
		3191 => "11111111",
		3192 => "11111111",
		3193 => "11111111",
		3194 => "11111111",
		3195 => "11111111",
		3196 => "11111111",
		3197 => "11111111",
		3198 => "11111111",
		3199 => "11111111",
		3200 => "11111111",
		3201 => "11111111",
		3202 => "11111111",
		3203 => "11111111",
		3204 => "11111111",
		3205 => "11111111",
		3206 => "11111111",
		3207 => "11111111",
		3208 => "11111111",
		3209 => "11111111",
		3210 => "11111111",
		3211 => "11111111",
		3212 => "11111111",
		3213 => "11111111",
		3214 => "11111111",
		3215 => "11111111",
		3216 => "11111111",
		3217 => "11111111",
		3218 => "11111111",
		3219 => "11111111",
		3220 => "11111111",
		3221 => "11111111",
		3222 => "11111111",
		3223 => "11111111",
		3224 => "11111111",
		3225 => "11111111",
		3226 => "11010001",
		3227 => "01001101",
		3228 => "01001101",
		3229 => "11010001",
		3230 => "11111111",
		3231 => "11111111",
		3232 => "11111111",
		3233 => "11100010",
		3234 => "01000111",
		3235 => "11000101",
		3236 => "11111111",
		3237 => "11111111",
		3238 => "11111111",
		3239 => "11111111",
		3240 => "11111111",
		3241 => "11111111",
		3242 => "11111111",
		3243 => "11111111",
		3244 => "11111111",
		3245 => "11111111",
		3246 => "11101110",
		3247 => "01001101",
		3248 => "01110000",
		3249 => "11000000",
		3250 => "11110011",
		3251 => "11111111",
		3252 => "11111111",
		3253 => "11111001",
		3254 => "10000111",
		3255 => "01010011",
		3256 => "01000111",
		3257 => "01000111",
		3258 => "01100100",
		3259 => "10101001",
		3260 => "11010001",
		3261 => "11111001",
		3262 => "11111111",
		3263 => "11111111",
		3264 => "11111111",
		3265 => "11111111",
		3266 => "11111111",
		3267 => "11111111",
		3268 => "11111111",
		3269 => "11111111",
		3270 => "11111111",
		3271 => "11111111",
		3272 => "11111111",
		3273 => "11111111",
		3274 => "11111111",
		3275 => "11111111",
		3276 => "11111111",
		3277 => "11111111",
		3278 => "11101110",
		3279 => "10011000",
		3280 => "01000111",
		3281 => "11011100",
		3282 => "11111111",
		3283 => "11111111",
		3284 => "11111111",
		3285 => "11111111",
		3286 => "11111111",
		3287 => "11111111",
		3288 => "11111111",
		3289 => "11111111",
		3290 => "11111111",
		3291 => "11111111",
		3292 => "11111111",
		3293 => "11000000",
		3294 => "11001011",
		3295 => "11111111",
		3296 => "11111111",
		3297 => "11111111",
		3298 => "11001011",
		3299 => "01000111",
		3300 => "10000111",
		3301 => "11111001",
		3302 => "11111111",
		3303 => "11111111",
		3304 => "11111111",
		3305 => "11111111",
		3306 => "11111111",
		3307 => "11111111",
		3308 => "11111111",
		3309 => "11101000",
		3310 => "01011110",
		3311 => "11110011",
		3312 => "11111111",
		3313 => "11111111",
		3314 => "11111111",
		3315 => "11111111",
		3316 => "11111111",
		3317 => "11111111",
		3318 => "11111111",
		3319 => "11111111",
		3320 => "11111111",
		3321 => "11111111",
		3322 => "11111111",
		3323 => "11111111",
		3324 => "11111111",
		3325 => "11111111",
		3326 => "11111111",
		3327 => "11111111",
		3328 => "11111111",
		3329 => "11111111",
		3330 => "11111111",
		3331 => "11111111",
		3332 => "11111111",
		3333 => "11111111",
		3334 => "11111111",
		3335 => "11111111",
		3336 => "11111111",
		3337 => "11111111",
		3338 => "11111111",
		3339 => "11111111",
		3340 => "11111111",
		3341 => "11111111",
		3342 => "11111111",
		3343 => "11111111",
		3344 => "11111111",
		3345 => "11111111",
		3346 => "11111111",
		3347 => "11111111",
		3348 => "11111111",
		3349 => "11111111",
		3350 => "11111111",
		3351 => "11111111",
		3352 => "11111111",
		3353 => "11111111",
		3354 => "11111111",
		3355 => "11000101",
		3356 => "01000111",
		3357 => "01010011",
		3358 => "11011100",
		3359 => "11111111",
		3360 => "11111111",
		3361 => "01100100",
		3362 => "11001011",
		3363 => "11111111",
		3364 => "11111111",
		3365 => "11111111",
		3366 => "11111111",
		3367 => "11111111",
		3368 => "11111111",
		3369 => "11111111",
		3370 => "11111111",
		3371 => "11111111",
		3372 => "11111111",
		3373 => "11111111",
		3374 => "10100011",
		3375 => "01001101",
		3376 => "11101110",
		3377 => "11111111",
		3378 => "11110011",
		3379 => "10111010",
		3380 => "10000001",
		3381 => "01001101",
		3382 => "01101010",
		3383 => "10101110",
		3384 => "10100011",
		3385 => "01011110",
		3386 => "01010011",
		3387 => "11101110",
		3388 => "11111111",
		3389 => "11111111",
		3390 => "11111111",
		3391 => "11111111",
		3392 => "11111111",
		3393 => "11111111",
		3394 => "11111111",
		3395 => "11111111",
		3396 => "11111111",
		3397 => "11111111",
		3398 => "11111111",
		3399 => "11111111",
		3400 => "11111111",
		3401 => "11111111",
		3402 => "11111111",
		3403 => "11111111",
		3404 => "11111111",
		3405 => "11111111",
		3406 => "11111111",
		3407 => "11110011",
		3408 => "01000111",
		3409 => "10101001",
		3410 => "11111111",
		3411 => "11111111",
		3412 => "11111111",
		3413 => "11111111",
		3414 => "11111111",
		3415 => "11111111",
		3416 => "11111111",
		3417 => "11111111",
		3418 => "11111111",
		3419 => "11111111",
		3420 => "11111111",
		3421 => "11111111",
		3422 => "01001101",
		3423 => "11011100",
		3424 => "11111111",
		3425 => "11101110",
		3426 => "01011110",
		3427 => "01000111",
		3428 => "10000001",
		3429 => "01111100",
		3430 => "11110011",
		3431 => "11111111",
		3432 => "11111111",
		3433 => "11111111",
		3434 => "11111111",
		3435 => "11111111",
		3436 => "11111111",
		3437 => "10011110",
		3438 => "01000111",
		3439 => "10001100",
		3440 => "11111111",
		3441 => "11111111",
		3442 => "11111111",
		3443 => "11111111",
		3444 => "11111111",
		3445 => "11111111",
		3446 => "11111111",
		3447 => "11111111",
		3448 => "11111111",
		3449 => "11111111",
		3450 => "11111111",
		3451 => "11111111",
		3452 => "11111111",
		3453 => "11111111",
		3454 => "11111111",
		3455 => "11111111",
		3456 => "11111111",
		3457 => "11111111",
		3458 => "11111111",
		3459 => "11111111",
		3460 => "11111111",
		3461 => "11111111",
		3462 => "11111111",
		3463 => "11111111",
		3464 => "11111111",
		3465 => "11111111",
		3466 => "11111111",
		3467 => "11111111",
		3468 => "11111111",
		3469 => "11111111",
		3470 => "11111111",
		3471 => "11111111",
		3472 => "11110011",
		3473 => "10101110",
		3474 => "10100011",
		3475 => "11000101",
		3476 => "11111111",
		3477 => "11111111",
		3478 => "11111111",
		3479 => "11111111",
		3480 => "11111111",
		3481 => "11111111",
		3482 => "11111111",
		3483 => "11111111",
		3484 => "10111010",
		3485 => "01000111",
		3486 => "01011110",
		3487 => "11101000",
		3488 => "11010001",
		3489 => "11011100",
		3490 => "11111111",
		3491 => "11111111",
		3492 => "11111111",
		3493 => "11111111",
		3494 => "11111111",
		3495 => "11111111",
		3496 => "11111111",
		3497 => "11111111",
		3498 => "11111111",
		3499 => "11111111",
		3500 => "11111111",
		3501 => "11111111",
		3502 => "11000000",
		3503 => "01000111",
		3504 => "11000101",
		3505 => "10001100",
		3506 => "01001101",
		3507 => "01000111",
		3508 => "01000111",
		3509 => "01000111",
		3510 => "11111111",
		3511 => "11111111",
		3512 => "11111111",
		3513 => "11010001",
		3514 => "01000111",
		3515 => "10111010",
		3516 => "11111111",
		3517 => "11111111",
		3518 => "11111111",
		3519 => "11101110",
		3520 => "11010001",
		3521 => "10111010",
		3522 => "10100011",
		3523 => "10000111",
		3524 => "01110101",
		3525 => "01110101",
		3526 => "01110101",
		3527 => "01110101",
		3528 => "01110101",
		3529 => "01110101",
		3530 => "01110101",
		3531 => "10000111",
		3532 => "10100011",
		3533 => "10100011",
		3534 => "11000000",
		3535 => "10000001",
		3536 => "01000111",
		3537 => "11010111",
		3538 => "11111111",
		3539 => "11111111",
		3540 => "11111111",
		3541 => "11111111",
		3542 => "11111111",
		3543 => "11111111",
		3544 => "11111111",
		3545 => "11111111",
		3546 => "11111111",
		3547 => "11111111",
		3548 => "11111111",
		3549 => "11111111",
		3550 => "11000000",
		3551 => "01011001",
		3552 => "10101001",
		3553 => "01110101",
		3554 => "01000111",
		3555 => "10011000",
		3556 => "11111111",
		3557 => "11111111",
		3558 => "11111111",
		3559 => "11111111",
		3560 => "11111111",
		3561 => "11111111",
		3562 => "11111111",
		3563 => "11100010",
		3564 => "01110000",
		3565 => "01010011",
		3566 => "01000111",
		3567 => "10011000",
		3568 => "11111111",
		3569 => "11111111",
		3570 => "11111111",
		3571 => "11111111",
		3572 => "11111111",
		3573 => "11111111",
		3574 => "11111111",
		3575 => "11111111",
		3576 => "11111111",
		3577 => "11111111",
		3578 => "11111111",
		3579 => "11111111",
		3580 => "11111111",
		3581 => "11111111",
		3582 => "11111111",
		3583 => "11111111",
		3584 => "11111111",
		3585 => "11111111",
		3586 => "11111111",
		3587 => "11111111",
		3588 => "11111111",
		3589 => "11111111",
		3590 => "11111111",
		3591 => "11111111",
		3592 => "11111111",
		3593 => "11111111",
		3594 => "11111111",
		3595 => "11111111",
		3596 => "11111111",
		3597 => "11111111",
		3598 => "11111111",
		3599 => "11101110",
		3600 => "01011110",
		3601 => "01000111",
		3602 => "01000111",
		3603 => "01000111",
		3604 => "10010011",
		3605 => "11111111",
		3606 => "11111111",
		3607 => "11111111",
		3608 => "11111111",
		3609 => "11111111",
		3610 => "11111111",
		3611 => "11111111",
		3612 => "11111111",
		3613 => "10100011",
		3614 => "01000111",
		3615 => "01011001",
		3616 => "01110000",
		3617 => "11111111",
		3618 => "11111111",
		3619 => "11111111",
		3620 => "11111111",
		3621 => "11111111",
		3622 => "11111111",
		3623 => "11111111",
		3624 => "11111111",
		3625 => "11111111",
		3626 => "11111111",
		3627 => "11111111",
		3628 => "11111111",
		3629 => "11111111",
		3630 => "11011100",
		3631 => "01000111",
		3632 => "01000111",
		3633 => "01010011",
		3634 => "10010011",
		3635 => "11101000",
		3636 => "11110011",
		3637 => "10011000",
		3638 => "11000000",
		3639 => "11111111",
		3640 => "11111111",
		3641 => "11101110",
		3642 => "01000111",
		3643 => "10001100",
		3644 => "10101001",
		3645 => "10000001",
		3646 => "01011110",
		3647 => "01000111",
		3648 => "01000111",
		3649 => "01000111",
		3650 => "01000111",
		3651 => "01011110",
		3652 => "01110101",
		3653 => "01110101",
		3654 => "01110101",
		3655 => "01110101",
		3656 => "01110101",
		3657 => "01110101",
		3658 => "01110101",
		3659 => "01110101",
		3660 => "01011110",
		3661 => "01000111",
		3662 => "01000111",
		3663 => "01000111",
		3664 => "10000001",
		3665 => "11111111",
		3666 => "11111111",
		3667 => "11111111",
		3668 => "11111111",
		3669 => "11111111",
		3670 => "11111111",
		3671 => "11111111",
		3672 => "11111111",
		3673 => "11111111",
		3674 => "11111111",
		3675 => "11111111",
		3676 => "11111111",
		3677 => "11111111",
		3678 => "11111111",
		3679 => "11101110",
		3680 => "10011000",
		3681 => "01001101",
		3682 => "01111100",
		3683 => "11111111",
		3684 => "11111111",
		3685 => "11111111",
		3686 => "11111111",
		3687 => "11111111",
		3688 => "11111111",
		3689 => "11111111",
		3690 => "10111010",
		3691 => "01010011",
		3692 => "10101001",
		3693 => "10010011",
		3694 => "01000111",
		3695 => "11010001",
		3696 => "11111111",
		3697 => "11111111",
		3698 => "11111111",
		3699 => "11111111",
		3700 => "11111111",
		3701 => "11111111",
		3702 => "11111111",
		3703 => "11111111",
		3704 => "11111111",
		3705 => "11111111",
		3706 => "11111111",
		3707 => "11111111",
		3708 => "11111111",
		3709 => "11111111",
		3710 => "11111111",
		3711 => "11111111",
		3712 => "11111111",
		3713 => "11111111",
		3714 => "11111111",
		3715 => "11111111",
		3716 => "11111111",
		3717 => "11111111",
		3718 => "11111111",
		3719 => "11111111",
		3720 => "11111111",
		3721 => "11111111",
		3722 => "11111111",
		3723 => "11111111",
		3724 => "11111111",
		3725 => "11111111",
		3726 => "11111001",
		3727 => "01110101",
		3728 => "10111010",
		3729 => "11111111",
		3730 => "11000101",
		3731 => "01010011",
		3732 => "01000111",
		3733 => "11011100",
		3734 => "11111111",
		3735 => "11111111",
		3736 => "11111111",
		3737 => "11111111",
		3738 => "11111111",
		3739 => "11111111",
		3740 => "11111111",
		3741 => "11111111",
		3742 => "01011110",
		3743 => "01111100",
		3744 => "11110011",
		3745 => "11111111",
		3746 => "11111111",
		3747 => "11111111",
		3748 => "11111111",
		3749 => "11111111",
		3750 => "11111111",
		3751 => "11111111",
		3752 => "11111111",
		3753 => "11111111",
		3754 => "11111111",
		3755 => "11111111",
		3756 => "11110011",
		3757 => "10011110",
		3758 => "01000111",
		3759 => "01000111",
		3760 => "01000111",
		3761 => "10101001",
		3762 => "11111111",
		3763 => "11111111",
		3764 => "11111111",
		3765 => "11111001",
		3766 => "10000001",
		3767 => "11111111",
		3768 => "11111111",
		3769 => "10100011",
		3770 => "01000111",
		3771 => "01000111",
		3772 => "01000111",
		3773 => "01011110",
		3774 => "10000111",
		3775 => "10101001",
		3776 => "11010001",
		3777 => "11100010",
		3778 => "11111111",
		3779 => "11111111",
		3780 => "11111111",
		3781 => "11111111",
		3782 => "11111111",
		3783 => "11111111",
		3784 => "11111111",
		3785 => "11111111",
		3786 => "11111111",
		3787 => "11111111",
		3788 => "11101110",
		3789 => "01011001",
		3790 => "01000111",
		3791 => "01000111",
		3792 => "01000111",
		3793 => "01101010",
		3794 => "11010001",
		3795 => "11111111",
		3796 => "11111111",
		3797 => "11111111",
		3798 => "11111111",
		3799 => "11111111",
		3800 => "11111111",
		3801 => "11111111",
		3802 => "11111111",
		3803 => "11111111",
		3804 => "11111111",
		3805 => "11111111",
		3806 => "11111111",
		3807 => "11111111",
		3808 => "11111111",
		3809 => "11101110",
		3810 => "11110011",
		3811 => "11111111",
		3812 => "11111111",
		3813 => "11111111",
		3814 => "11111111",
		3815 => "11111111",
		3816 => "11110011",
		3817 => "10000001",
		3818 => "01100100",
		3819 => "11010111",
		3820 => "11111111",
		3821 => "01011001",
		3822 => "01010011",
		3823 => "11111111",
		3824 => "11111111",
		3825 => "11111111",
		3826 => "11111111",
		3827 => "11111111",
		3828 => "11111111",
		3829 => "11111111",
		3830 => "11111111",
		3831 => "11111111",
		3832 => "11111111",
		3833 => "11111111",
		3834 => "11111111",
		3835 => "11111111",
		3836 => "11111111",
		3837 => "11111111",
		3838 => "11111111",
		3839 => "11111111",
		3840 => "11111111",
		3841 => "11111111",
		3842 => "11111111",
		3843 => "11111111",
		3844 => "11111111",
		3845 => "11111111",
		3846 => "11111111",
		3847 => "11111111",
		3848 => "11111111",
		3849 => "11111111",
		3850 => "11111111",
		3851 => "11111111",
		3852 => "11111111",
		3853 => "11111111",
		3854 => "10011000",
		3855 => "10111010",
		3856 => "11111111",
		3857 => "11111111",
		3858 => "11111111",
		3859 => "11010111",
		3860 => "01000111",
		3861 => "10111010",
		3862 => "11111111",
		3863 => "11111111",
		3864 => "11111111",
		3865 => "11111111",
		3866 => "11111111",
		3867 => "11111111",
		3868 => "11111111",
		3869 => "11000101",
		3870 => "10010011",
		3871 => "11111111",
		3872 => "11111111",
		3873 => "11111111",
		3874 => "11111111",
		3875 => "11111111",
		3876 => "11111111",
		3877 => "11111111",
		3878 => "11111111",
		3879 => "11111111",
		3880 => "11111111",
		3881 => "11111111",
		3882 => "11111111",
		3883 => "11001011",
		3884 => "01011001",
		3885 => "01000111",
		3886 => "10001100",
		3887 => "10110100",
		3888 => "01110101",
		3889 => "01000111",
		3890 => "10111010",
		3891 => "11111111",
		3892 => "11111111",
		3893 => "11111111",
		3894 => "01110101",
		3895 => "11111111",
		3896 => "11111111",
		3897 => "10010011",
		3898 => "01000111",
		3899 => "01000111",
		3900 => "10011000",
		3901 => "11111111",
		3902 => "11111111",
		3903 => "11111111",
		3904 => "11111111",
		3905 => "11111111",
		3906 => "11111111",
		3907 => "11111111",
		3908 => "11111111",
		3909 => "11111111",
		3910 => "11111111",
		3911 => "11111111",
		3912 => "11111111",
		3913 => "11111001",
		3914 => "11010001",
		3915 => "11101110",
		3916 => "11101000",
		3917 => "01010011",
		3918 => "01000111",
		3919 => "01000111",
		3920 => "01110000",
		3921 => "01011001",
		3922 => "01000111",
		3923 => "01111100",
		3924 => "11110011",
		3925 => "11111111",
		3926 => "11111111",
		3927 => "11111111",
		3928 => "11111111",
		3929 => "11111111",
		3930 => "11111111",
		3931 => "11111111",
		3932 => "11111111",
		3933 => "11111111",
		3934 => "11111111",
		3935 => "11111111",
		3936 => "11111111",
		3937 => "11111111",
		3938 => "11111111",
		3939 => "11111111",
		3940 => "11111111",
		3941 => "11111111",
		3942 => "11111111",
		3943 => "11010001",
		3944 => "01011001",
		3945 => "10010011",
		3946 => "11111001",
		3947 => "11111111",
		3948 => "11010001",
		3949 => "01000111",
		3950 => "10001100",
		3951 => "11111111",
		3952 => "11111111",
		3953 => "11111111",
		3954 => "11111111",
		3955 => "11111111",
		3956 => "11111111",
		3957 => "11111111",
		3958 => "11111111",
		3959 => "11111111",
		3960 => "11111111",
		3961 => "11111111",
		3962 => "11111111",
		3963 => "11111111",
		3964 => "11111111",
		3965 => "11111111",
		3966 => "11111111",
		3967 => "11111111",
		3968 => "11111111",
		3969 => "11111111",
		3970 => "11111111",
		3971 => "11111111",
		3972 => "11111111",
		3973 => "11111111",
		3974 => "11111111",
		3975 => "11111111",
		3976 => "11111111",
		3977 => "11111111",
		3978 => "11111111",
		3979 => "11111111",
		3980 => "11111111",
		3981 => "11000101",
		3982 => "01000111",
		3983 => "10011110",
		3984 => "11111001",
		3985 => "11111111",
		3986 => "11111111",
		3987 => "11111111",
		3988 => "01011110",
		3989 => "11011100",
		3990 => "11111111",
		3991 => "11111111",
		3992 => "11111111",
		3993 => "11111111",
		3994 => "11111111",
		3995 => "11111001",
		3996 => "10110100",
		3997 => "11110100",
		3998 => "11111111",
		3999 => "11111111",
		4000 => "11111111",
		4001 => "11111111",
		4002 => "11111111",
		4003 => "11111111",
		4004 => "11111111",
		4005 => "11111111",
		4006 => "11111111",
		4007 => "11111111",
		4008 => "11111111",
		4009 => "11111111",
		4010 => "10101110",
		4011 => "01000111",
		4012 => "01100100",
		4013 => "11010111",
		4014 => "11111111",
		4015 => "11111111",
		4016 => "11111001",
		4017 => "01011001",
		4018 => "01100100",
		4019 => "11111111",
		4020 => "11111111",
		4021 => "11101110",
		4022 => "01000111",
		4023 => "01110101",
		4024 => "11010111",
		4025 => "11111111",
		4026 => "11111001",
		4027 => "10001100",
		4028 => "01000111",
		4029 => "11101000",
		4030 => "11111111",
		4031 => "11111111",
		4032 => "11100010",
		4033 => "11000101",
		4034 => "10100011",
		4035 => "01111100",
		4036 => "01011110",
		4037 => "01000111",
		4038 => "01000111",
		4039 => "01000111",
		4040 => "01000111",
		4041 => "01000111",
		4042 => "01000111",
		4043 => "01000111",
		4044 => "01000111",
		4045 => "01000111",
		4046 => "01011110",
		4047 => "11101110",
		4048 => "11111111",
		4049 => "11111111",
		4050 => "10101001",
		4051 => "01001101",
		4052 => "01011001",
		4053 => "11010001",
		4054 => "11111111",
		4055 => "11111111",
		4056 => "11111111",
		4057 => "11111111",
		4058 => "11111111",
		4059 => "11111111",
		4060 => "11111111",
		4061 => "11111111",
		4062 => "11111111",
		4063 => "11111111",
		4064 => "11111111",
		4065 => "11111111",
		4066 => "11111111",
		4067 => "11110011",
		4068 => "10011110",
		4069 => "11110011",
		4070 => "10011110",
		4071 => "01011001",
		4072 => "11001011",
		4073 => "11111111",
		4074 => "11111111",
		4075 => "11111111",
		4076 => "10011110",
		4077 => "01000111",
		4078 => "11000000",
		4079 => "11111111",
		4080 => "11111111",
		4081 => "11111111",
		4082 => "11000000",
		4083 => "11111111",
		4084 => "11111111",
		4085 => "11111111",
		4086 => "11111111",
		4087 => "11111111",
		4088 => "11111111",
		4089 => "11111111",
		4090 => "11111111",
		4091 => "11111111",
		4092 => "11111111",
		4093 => "11111111",
		4094 => "11111111",
		4095 => "11111111",
		4096 => "11111111",
		4097 => "11111111",
		4098 => "11111111",
		4099 => "11111111",
		4100 => "11111111",
		4101 => "11111111",
		4102 => "11111111",
		4103 => "11111111",
		4104 => "11111111",
		4105 => "11111111",
		4106 => "11111111",
		4107 => "11111111",
		4108 => "11111111",
		4109 => "01010011",
		4110 => "01011001",
		4111 => "01000111",
		4112 => "01110000",
		4113 => "11100010",
		4114 => "11111111",
		4115 => "11111001",
		4116 => "01010011",
		4117 => "01110101",
		4118 => "01110101",
		4119 => "01110101",
		4120 => "01110101",
		4121 => "01110101",
		4122 => "01110101",
		4123 => "01011110",
		4124 => "10011000",
		4125 => "11111111",
		4126 => "11111111",
		4127 => "11111111",
		4128 => "11111111",
		4129 => "11111111",
		4130 => "11111111",
		4131 => "11111111",
		4132 => "11111111",
		4133 => "11111111",
		4134 => "11111111",
		4135 => "11111111",
		4136 => "11111111",
		4137 => "10010011",
		4138 => "01000111",
		4139 => "10001100",
		4140 => "11111001",
		4141 => "11111111",
		4142 => "11111111",
		4143 => "11111111",
		4144 => "11111111",
		4145 => "10011000",
		4146 => "01000111",
		4147 => "11111111",
		4148 => "11111111",
		4149 => "11111001",
		4150 => "10100011",
		4151 => "01011110",
		4152 => "01010011",
		4153 => "11110011",
		4154 => "11111111",
		4155 => "11000101",
		4156 => "01000111",
		4157 => "10001100",
		4158 => "01111100",
		4159 => "01010011",
		4160 => "01000111",
		4161 => "01000111",
		4162 => "01000111",
		4163 => "01100100",
		4164 => "10000111",
		4165 => "10100011",
		4166 => "10100011",
		4167 => "10100011",
		4168 => "11001011",
		4169 => "11010001",
		4170 => "01000111",
		4171 => "01111100",
		4172 => "10011000",
		4173 => "01000111",
		4174 => "10011110",
		4175 => "11111111",
		4176 => "11111111",
		4177 => "11111111",
		4178 => "11111111",
		4179 => "11100010",
		4180 => "01101010",
		4181 => "01001101",
		4182 => "10111010",
		4183 => "11111111",
		4184 => "11111111",
		4185 => "11111111",
		4186 => "11111111",
		4187 => "11111111",
		4188 => "11111111",
		4189 => "11111111",
		4190 => "11111111",
		4191 => "11111111",
		4192 => "11111111",
		4193 => "11111111",
		4194 => "11111111",
		4195 => "11111111",
		4196 => "10100011",
		4197 => "01000111",
		4198 => "01111100",
		4199 => "11101110",
		4200 => "11111111",
		4201 => "11111111",
		4202 => "11111111",
		4203 => "11111111",
		4204 => "01011110",
		4205 => "01001101",
		4206 => "11111001",
		4207 => "11111111",
		4208 => "11111111",
		4209 => "11111111",
		4210 => "11100010",
		4211 => "11101000",
		4212 => "11111111",
		4213 => "11111111",
		4214 => "11111111",
		4215 => "11111111",
		4216 => "11111111",
		4217 => "11111111",
		4218 => "11111111",
		4219 => "11111111",
		4220 => "11111111",
		4221 => "11111111",
		4222 => "11111111",
		4223 => "11111111",
		4224 => "11111111",
		4225 => "11111111",
		4226 => "11111111",
		4227 => "11111111",
		4228 => "11111111",
		4229 => "11111111",
		4230 => "11111111",
		4231 => "11111111",
		4232 => "11111111",
		4233 => "11111111",
		4234 => "11111111",
		4235 => "11111111",
		4236 => "11111111",
		4237 => "11111111",
		4238 => "11111111",
		4239 => "11111111",
		4240 => "10111010",
		4241 => "01010011",
		4242 => "01000111",
		4243 => "01010011",
		4244 => "11110011",
		4245 => "11111111",
		4246 => "11111111",
		4247 => "11111111",
		4248 => "11111111",
		4249 => "11111111",
		4250 => "11111111",
		4251 => "11111111",
		4252 => "11111111",
		4253 => "11111111",
		4254 => "11111111",
		4255 => "11111111",
		4256 => "11111111",
		4257 => "11111111",
		4258 => "11111111",
		4259 => "11111111",
		4260 => "11111111",
		4261 => "11111111",
		4262 => "11111111",
		4263 => "11011100",
		4264 => "01000111",
		4265 => "10001100",
		4266 => "11111111",
		4267 => "11111111",
		4268 => "11111111",
		4269 => "11111111",
		4270 => "11111111",
		4271 => "11111111",
		4272 => "11111111",
		4273 => "10101110",
		4274 => "10010011",
		4275 => "10011110",
		4276 => "01011110",
		4277 => "01001101",
		4278 => "11111111",
		4279 => "10011110",
		4280 => "01000111",
		4281 => "01110000",
		4282 => "11000101",
		4283 => "10101001",
		4284 => "01110101",
		4285 => "01000111",
		4286 => "10011000",
		4287 => "11111111",
		4288 => "11111111",
		4289 => "11111001",
		4290 => "11001011",
		4291 => "10100011",
		4292 => "10000111",
		4293 => "01110101",
		4294 => "01000111",
		4295 => "01000111",
		4296 => "01000111",
		4297 => "01000111",
		4298 => "01000111",
		4299 => "01000111",
		4300 => "01110000",
		4301 => "01100100",
		4302 => "01011110",
		4303 => "11111111",
		4304 => "11111111",
		4305 => "11111111",
		4306 => "11111111",
		4307 => "11111111",
		4308 => "11111111",
		4309 => "11111001",
		4310 => "01101010",
		4311 => "01010011",
		4312 => "11101110",
		4313 => "11111111",
		4314 => "11111111",
		4315 => "11111111",
		4316 => "11111111",
		4317 => "11111111",
		4318 => "11111111",
		4319 => "11111111",
		4320 => "11111111",
		4321 => "11111111",
		4322 => "11111111",
		4323 => "11111111",
		4324 => "11111111",
		4325 => "11101110",
		4326 => "10111010",
		4327 => "11111111",
		4328 => "11111111",
		4329 => "11111111",
		4330 => "11111111",
		4331 => "10100011",
		4332 => "01000111",
		4333 => "10110100",
		4334 => "11111111",
		4335 => "11111111",
		4336 => "10101110",
		4337 => "01010011",
		4338 => "10101001",
		4339 => "11010001",
		4340 => "11100010",
		4341 => "11111111",
		4342 => "11111111",
		4343 => "11111111",
		4344 => "11111111",
		4345 => "11111111",
		4346 => "11111111",
		4347 => "11111111",
		4348 => "11111111",
		4349 => "11111111",
		4350 => "11111111",
		4351 => "11111111",
		4352 => "11111111",
		4353 => "11111111",
		4354 => "11111111",
		4355 => "11111111",
		4356 => "11111111",
		4357 => "11111111",
		4358 => "11111111",
		4359 => "11111111",
		4360 => "11111111",
		4361 => "11111111",
		4362 => "11111111",
		4363 => "11111111",
		4364 => "11111111",
		4365 => "11111111",
		4366 => "11111111",
		4367 => "11111111",
		4368 => "11111111",
		4369 => "11100010",
		4370 => "01110000",
		4371 => "01000111",
		4372 => "01011001",
		4373 => "11001011",
		4374 => "11111111",
		4375 => "11111111",
		4376 => "11111111",
		4377 => "11111111",
		4378 => "11111111",
		4379 => "11111111",
		4380 => "11111111",
		4381 => "11111111",
		4382 => "11111111",
		4383 => "11111111",
		4384 => "11111111",
		4385 => "11111111",
		4386 => "11111111",
		4387 => "11111111",
		4388 => "11111111",
		4389 => "11111111",
		4390 => "11111111",
		4391 => "10000001",
		4392 => "01010011",
		4393 => "11111001",
		4394 => "11111111",
		4395 => "11111111",
		4396 => "11111111",
		4397 => "11111111",
		4398 => "11111111",
		4399 => "11111111",
		4400 => "11111111",
		4401 => "11111111",
		4402 => "11111111",
		4403 => "11111111",
		4404 => "11011100",
		4405 => "01000111",
		4406 => "11111111",
		4407 => "10110100",
		4408 => "01110101",
		4409 => "01100100",
		4410 => "01000111",
		4411 => "11000101",
		4412 => "11111111",
		4413 => "10010011",
		4414 => "01001101",
		4415 => "10011110",
		4416 => "01110000",
		4417 => "01000111",
		4418 => "01000111",
		4419 => "01000111",
		4420 => "01010011",
		4421 => "01000111",
		4422 => "01000111",
		4423 => "01000111",
		4424 => "10000001",
		4425 => "11010001",
		4426 => "01000111",
		4427 => "11000101",
		4428 => "11111111",
		4429 => "11111111",
		4430 => "11111111",
		4431 => "11111111",
		4432 => "11111111",
		4433 => "11111111",
		4434 => "11111111",
		4435 => "11111111",
		4436 => "11111111",
		4437 => "11111111",
		4438 => "11100010",
		4439 => "01001101",
		4440 => "10011000",
		4441 => "11111111",
		4442 => "11111111",
		4443 => "11111111",
		4444 => "11111111",
		4445 => "11111111",
		4446 => "11111111",
		4447 => "11111111",
		4448 => "11111111",
		4449 => "11111111",
		4450 => "11111111",
		4451 => "11111111",
		4452 => "11111111",
		4453 => "11111111",
		4454 => "11111111",
		4455 => "11111111",
		4456 => "11111111",
		4457 => "11111111",
		4458 => "11111111",
		4459 => "01100100",
		4460 => "01000111",
		4461 => "11101110",
		4462 => "11101110",
		4463 => "01111100",
		4464 => "01101010",
		4465 => "11100010",
		4466 => "11111111",
		4467 => "11111111",
		4468 => "11111111",
		4469 => "11111111",
		4470 => "11111111",
		4471 => "11111111",
		4472 => "11111111",
		4473 => "11111111",
		4474 => "11111111",
		4475 => "11111111",
		4476 => "11111111",
		4477 => "11111111",
		4478 => "11111111",
		4479 => "11111111",
		4480 => "11111111",
		4481 => "11111111",
		4482 => "11111111",
		4483 => "11111111",
		4484 => "11111111",
		4485 => "11111111",
		4486 => "11111111",
		4487 => "11111111",
		4488 => "11111111",
		4489 => "11111111",
		4490 => "11111111",
		4491 => "11111111",
		4492 => "11111111",
		4493 => "11111111",
		4494 => "11111111",
		4495 => "11111111",
		4496 => "11111111",
		4497 => "11111111",
		4498 => "11111111",
		4499 => "10101001",
		4500 => "01000111",
		4501 => "01000111",
		4502 => "10010011",
		4503 => "11111001",
		4504 => "11010001",
		4505 => "11010111",
		4506 => "11111111",
		4507 => "11111111",
		4508 => "11111111",
		4509 => "11111111",
		4510 => "11111111",
		4511 => "11111111",
		4512 => "11111111",
		4513 => "11111111",
		4514 => "11111111",
		4515 => "11111111",
		4516 => "11111111",
		4517 => "11111111",
		4518 => "11111111",
		4519 => "01000111",
		4520 => "10000111",
		4521 => "11111111",
		4522 => "11111111",
		4523 => "11111111",
		4524 => "11111111",
		4525 => "11111111",
		4526 => "11111111",
		4527 => "11111111",
		4528 => "11111111",
		4529 => "11111111",
		4530 => "11111111",
		4531 => "11111111",
		4532 => "11111111",
		4533 => "01011001",
		4534 => "01110101",
		4535 => "10011000",
		4536 => "11110011",
		4537 => "11111001",
		4538 => "01011001",
		4539 => "01110000",
		4540 => "10101110",
		4541 => "01011110",
		4542 => "01000111",
		4543 => "01000111",
		4544 => "01000111",
		4545 => "01000111",
		4546 => "01100100",
		4547 => "11101000",
		4548 => "10000111",
		4549 => "01011001",
		4550 => "11101110",
		4551 => "11111111",
		4552 => "11010111",
		4553 => "10100011",
		4554 => "01011001",
		4555 => "11111111",
		4556 => "11111111",
		4557 => "11111111",
		4558 => "11111111",
		4559 => "11111111",
		4560 => "11111111",
		4561 => "11111111",
		4562 => "11111111",
		4563 => "11111111",
		4564 => "11111111",
		4565 => "11111111",
		4566 => "11111111",
		4567 => "01110101",
		4568 => "01100100",
		4569 => "11111111",
		4570 => "11111111",
		4571 => "11111111",
		4572 => "11111111",
		4573 => "11111111",
		4574 => "11111111",
		4575 => "11111111",
		4576 => "11111111",
		4577 => "11111111",
		4578 => "11111111",
		4579 => "11111111",
		4580 => "11111111",
		4581 => "11111111",
		4582 => "11111111",
		4583 => "11111111",
		4584 => "11111111",
		4585 => "11111111",
		4586 => "11100010",
		4587 => "01000111",
		4588 => "01110000",
		4589 => "11001011",
		4590 => "01011001",
		4591 => "10011110",
		4592 => "11111001",
		4593 => "11111111",
		4594 => "11111111",
		4595 => "11111111",
		4596 => "11111111",
		4597 => "11111111",
		4598 => "11111111",
		4599 => "11111111",
		4600 => "11111111",
		4601 => "11111111",
		4602 => "11111111",
		4603 => "11111111",
		4604 => "11111111",
		4605 => "11111111",
		4606 => "11111111",
		4607 => "11111111",
		4608 => "11111111",
		4609 => "11111111",
		4610 => "11111111",
		4611 => "11111111",
		4612 => "11111111",
		4613 => "11111111",
		4614 => "11111111",
		4615 => "11111111",
		4616 => "11111111",
		4617 => "11111111",
		4618 => "11111111",
		4619 => "11111111",
		4620 => "11111111",
		4621 => "11111111",
		4622 => "11111111",
		4623 => "11111111",
		4624 => "11111111",
		4625 => "11111111",
		4626 => "11111111",
		4627 => "11111111",
		4628 => "11010111",
		4629 => "01100100",
		4630 => "01000111",
		4631 => "01011001",
		4632 => "01100100",
		4633 => "11111001",
		4634 => "11111111",
		4635 => "11111111",
		4636 => "11111111",
		4637 => "11111111",
		4638 => "11111111",
		4639 => "11111111",
		4640 => "11111111",
		4641 => "11111111",
		4642 => "11111111",
		4643 => "11101000",
		4644 => "11010001",
		4645 => "11010001",
		4646 => "11011100",
		4647 => "01001101",
		4648 => "10000111",
		4649 => "11111111",
		4650 => "11111111",
		4651 => "11111111",
		4652 => "11111111",
		4653 => "11111111",
		4654 => "11111111",
		4655 => "11111111",
		4656 => "11111111",
		4657 => "11111111",
		4658 => "11111111",
		4659 => "11111111",
		4660 => "11101110",
		4661 => "01000111",
		4662 => "01011110",
		4663 => "01000111",
		4664 => "01011110",
		4665 => "11101110",
		4666 => "01100100",
		4667 => "01000111",
		4668 => "01000111",
		4669 => "10000001",
		4670 => "11000000",
		4671 => "11101000",
		4672 => "10111010",
		4673 => "10000001",
		4674 => "01000111",
		4675 => "01000111",
		4676 => "01000111",
		4677 => "01110000",
		4678 => "11111111",
		4679 => "10101110",
		4680 => "01000111",
		4681 => "01000111",
		4682 => "01000111",
		4683 => "11111001",
		4684 => "11111111",
		4685 => "11111111",
		4686 => "11111111",
		4687 => "11111111",
		4688 => "11111111",
		4689 => "11111111",
		4690 => "11111111",
		4691 => "11111111",
		4692 => "11111111",
		4693 => "11111111",
		4694 => "11111111",
		4695 => "10000111",
		4696 => "01011110",
		4697 => "11111111",
		4698 => "11010001",
		4699 => "10100011",
		4700 => "10101001",
		4701 => "11010111",
		4702 => "11111111",
		4703 => "11111111",
		4704 => "11111111",
		4705 => "11111111",
		4706 => "11111111",
		4707 => "11111111",
		4708 => "11111111",
		4709 => "11111111",
		4710 => "11111111",
		4711 => "11111111",
		4712 => "11111111",
		4713 => "11111111",
		4714 => "10101001",
		4715 => "01000111",
		4716 => "01011001",
		4717 => "01011001",
		4718 => "11010001",
		4719 => "11111111",
		4720 => "11111111",
		4721 => "11111111",
		4722 => "11111111",
		4723 => "11111111",
		4724 => "11111111",
		4725 => "11111111",
		4726 => "11111001",
		4727 => "11111111",
		4728 => "11111111",
		4729 => "11111111",
		4730 => "11111111",
		4731 => "11111111",
		4732 => "11111111",
		4733 => "11111111",
		4734 => "11111111",
		4735 => "11111111",
		4736 => "11111111",
		4737 => "11111111",
		4738 => "11111111",
		4739 => "11111111",
		4740 => "11111111",
		4741 => "11111111",
		4742 => "11111111",
		4743 => "11111111",
		4744 => "11111111",
		4745 => "11111111",
		4746 => "11111111",
		4747 => "10011110",
		4748 => "01010011",
		4749 => "10000001",
		4750 => "11101110",
		4751 => "11111111",
		4752 => "11111111",
		4753 => "11111111",
		4754 => "11111111",
		4755 => "11111111",
		4756 => "11111111",
		4757 => "11111001",
		4758 => "10000001",
		4759 => "01001101",
		4760 => "11100010",
		4761 => "11111111",
		4762 => "11111111",
		4763 => "11111111",
		4764 => "11111111",
		4765 => "11111111",
		4766 => "11111111",
		4767 => "11111111",
		4768 => "11111111",
		4769 => "11001011",
		4770 => "01111100",
		4771 => "01000111",
		4772 => "01000111",
		4773 => "01000111",
		4774 => "01000111",
		4775 => "01000111",
		4776 => "01000111",
		4777 => "11001011",
		4778 => "11111111",
		4779 => "11111111",
		4780 => "11111111",
		4781 => "11111111",
		4782 => "11111111",
		4783 => "11111111",
		4784 => "11111111",
		4785 => "11111111",
		4786 => "11111111",
		4787 => "11111111",
		4788 => "11111111",
		4789 => "11010001",
		4790 => "11111111",
		4791 => "11000000",
		4792 => "01000111",
		4793 => "01000111",
		4794 => "01000111",
		4795 => "10001100",
		4796 => "11011100",
		4797 => "11111111",
		4798 => "11111111",
		4799 => "11111111",
		4800 => "11111111",
		4801 => "11111111",
		4802 => "11101110",
		4803 => "10011110",
		4804 => "01010011",
		4805 => "01000111",
		4806 => "10001100",
		4807 => "01001101",
		4808 => "01111100",
		4809 => "11101000",
		4810 => "10101001",
		4811 => "11111111",
		4812 => "11111111",
		4813 => "11111111",
		4814 => "11111111",
		4815 => "11111111",
		4816 => "11111111",
		4817 => "11111111",
		4818 => "11111111",
		4819 => "11111111",
		4820 => "11111111",
		4821 => "11111111",
		4822 => "11010111",
		4823 => "01000111",
		4824 => "01001101",
		4825 => "01000111",
		4826 => "01000111",
		4827 => "01000111",
		4828 => "01000111",
		4829 => "01000111",
		4830 => "10101001",
		4831 => "11111001",
		4832 => "11111111",
		4833 => "11111111",
		4834 => "11111111",
		4835 => "11111111",
		4836 => "11111111",
		4837 => "11111111",
		4838 => "11111111",
		4839 => "11111111",
		4840 => "11111111",
		4841 => "11111111",
		4842 => "01110000",
		4843 => "01000111",
		4844 => "10000111",
		4845 => "11110011",
		4846 => "11111111",
		4847 => "11111111",
		4848 => "11111111",
		4849 => "11111111",
		4850 => "11111111",
		4851 => "11111111",
		4852 => "11111111",
		4853 => "11010001",
		4854 => "10101110",
		4855 => "11111111",
		4856 => "11111111",
		4857 => "11111111",
		4858 => "11111111",
		4859 => "11111111",
		4860 => "11111111",
		4861 => "11111111",
		4862 => "11111111",
		4863 => "11111111",
		4864 => "11111111",
		4865 => "11111111",
		4866 => "11111111",
		4867 => "11111111",
		4868 => "11111111",
		4869 => "11111111",
		4870 => "11111111",
		4871 => "11111111",
		4872 => "11111111",
		4873 => "11111111",
		4874 => "10001100",
		4875 => "01011110",
		4876 => "01101010",
		4877 => "01000111",
		4878 => "01011001",
		4879 => "11101110",
		4880 => "11111111",
		4881 => "11111111",
		4882 => "11111111",
		4883 => "11111111",
		4884 => "11111111",
		4885 => "11111111",
		4886 => "10010011",
		4887 => "10111010",
		4888 => "11111111",
		4889 => "11111111",
		4890 => "11111111",
		4891 => "11111111",
		4892 => "11111111",
		4893 => "11111111",
		4894 => "11111111",
		4895 => "11111111",
		4896 => "11111001",
		4897 => "01000111",
		4898 => "01011001",
		4899 => "10100011",
		4900 => "11010001",
		4901 => "11010001",
		4902 => "10111010",
		4903 => "01110101",
		4904 => "01000111",
		4905 => "01000111",
		4906 => "01101010",
		4907 => "01110101",
		4908 => "01110101",
		4909 => "01110101",
		4910 => "01110101",
		4911 => "01110101",
		4912 => "10011110",
		4913 => "11010001",
		4914 => "11111111",
		4915 => "11111111",
		4916 => "11111111",
		4917 => "11111111",
		4918 => "11111111",
		4919 => "11111111",
		4920 => "01000111",
		4921 => "01100100",
		4922 => "11010111",
		4923 => "11111111",
		4924 => "10111010",
		4925 => "10011000",
		4926 => "10001100",
		4927 => "11001011",
		4928 => "11111111",
		4929 => "11111111",
		4930 => "11111111",
		4931 => "11011100",
		4932 => "11000101",
		4933 => "10011000",
		4934 => "01000111",
		4935 => "01000111",
		4936 => "11010111",
		4937 => "11111111",
		4938 => "11111111",
		4939 => "11111111",
		4940 => "11111111",
		4941 => "11111111",
		4942 => "11111111",
		4943 => "11000101",
		4944 => "10100011",
		4945 => "10100011",
		4946 => "10100011",
		4947 => "10100011",
		4948 => "10100011",
		4949 => "10100011",
		4950 => "01011001",
		4951 => "01000111",
		4952 => "01001101",
		4953 => "10001100",
		4954 => "11100010",
		4955 => "11111111",
		4956 => "11101110",
		4957 => "11000000",
		4958 => "01000111",
		4959 => "01101010",
		4960 => "11100010",
		4961 => "11111111",
		4962 => "11111111",
		4963 => "11111111",
		4964 => "11111111",
		4965 => "11111111",
		4966 => "11111111",
		4967 => "11111111",
		4968 => "11111111",
		4969 => "11101000",
		4970 => "01010011",
		4971 => "10111010",
		4972 => "11111111",
		4973 => "11111111",
		4974 => "11111111",
		4975 => "11111111",
		4976 => "11111111",
		4977 => "11111111",
		4978 => "11111111",
		4979 => "11111111",
		4980 => "11111111",
		4981 => "11000000",
		4982 => "01011001",
		4983 => "11111001",
		4984 => "11111111",
		4985 => "11111111",
		4986 => "11111111",
		4987 => "11111111",
		4988 => "11111111",
		4989 => "11111111",
		4990 => "11111111",
		4991 => "11111111",
		4992 => "11111111",
		4993 => "11111111",
		4994 => "11111111",
		4995 => "11111111",
		4996 => "11111111",
		4997 => "11111111",
		4998 => "11111111",
		4999 => "11111111",
		5000 => "11111111",
		5001 => "11010111",
		5002 => "01111100",
		5003 => "11111001",
		5004 => "11111111",
		5005 => "10011000",
		5006 => "01000111",
		5007 => "10011110",
		5008 => "11111111",
		5009 => "11111111",
		5010 => "11111111",
		5011 => "11111111",
		5012 => "11111111",
		5013 => "11111111",
		5014 => "11001011",
		5015 => "11111111",
		5016 => "11111111",
		5017 => "11111111",
		5018 => "11111111",
		5019 => "11111111",
		5020 => "11111111",
		5021 => "11111111",
		5022 => "11111111",
		5023 => "11101000",
		5024 => "01100100",
		5025 => "10101001",
		5026 => "11111111",
		5027 => "11111111",
		5028 => "11111111",
		5029 => "11111111",
		5030 => "11111111",
		5031 => "11111111",
		5032 => "11010001",
		5033 => "01010011",
		5034 => "01000111",
		5035 => "01100100",
		5036 => "01110101",
		5037 => "01110101",
		5038 => "01110101",
		5039 => "01011110",
		5040 => "01000111",
		5041 => "01000111",
		5042 => "01101010",
		5043 => "11101000",
		5044 => "11111111",
		5045 => "11111111",
		5046 => "11111111",
		5047 => "11000000",
		5048 => "01000111",
		5049 => "11000000",
		5050 => "11110011",
		5051 => "01110000",
		5052 => "01000111",
		5053 => "01011110",
		5054 => "01000111",
		5055 => "01000111",
		5056 => "10011110",
		5057 => "10011000",
		5058 => "01001101",
		5059 => "01000111",
		5060 => "01000111",
		5061 => "01010011",
		5062 => "01110000",
		5063 => "01000111",
		5064 => "11000000",
		5065 => "11111111",
		5066 => "11111111",
		5067 => "11111111",
		5068 => "11111001",
		5069 => "10100011",
		5070 => "01010011",
		5071 => "01000111",
		5072 => "01000111",
		5073 => "01000111",
		5074 => "01000111",
		5075 => "01000111",
		5076 => "01000111",
		5077 => "01000111",
		5078 => "01000111",
		5079 => "01011001",
		5080 => "11011100",
		5081 => "11111111",
		5082 => "11111111",
		5083 => "11111111",
		5084 => "11111111",
		5085 => "11111111",
		5086 => "11010001",
		5087 => "01010011",
		5088 => "01001101",
		5089 => "11001011",
		5090 => "11111111",
		5091 => "11111111",
		5092 => "11111111",
		5093 => "11111111",
		5094 => "11111111",
		5095 => "11111111",
		5096 => "11111111",
		5097 => "11111001",
		5098 => "11101110",
		5099 => "11111111",
		5100 => "11111111",
		5101 => "11111111",
		5102 => "11111111",
		5103 => "11111111",
		5104 => "11111111",
		5105 => "11111111",
		5106 => "11111111",
		5107 => "11000101",
		5108 => "01110101",
		5109 => "01000111",
		5110 => "01000111",
		5111 => "10111010",
		5112 => "11111111",
		5113 => "11111111",
		5114 => "11111111",
		5115 => "11111111",
		5116 => "11111111",
		5117 => "11111111",
		5118 => "11111111",
		5119 => "11111111",
		5120 => "11111111",
		5121 => "11111111",
		5122 => "11111111",
		5123 => "11111111",
		5124 => "11111111",
		5125 => "11111111",
		5126 => "11111111",
		5127 => "11111111",
		5128 => "11111111",
		5129 => "01111100",
		5130 => "11101110",
		5131 => "11111111",
		5132 => "11111111",
		5133 => "11111111",
		5134 => "10011000",
		5135 => "10001100",
		5136 => "11111111",
		5137 => "11111111",
		5138 => "11111111",
		5139 => "11111111",
		5140 => "11111111",
		5141 => "11111111",
		5142 => "11111111",
		5143 => "11111111",
		5144 => "11111111",
		5145 => "11111111",
		5146 => "11111111",
		5147 => "11111111",
		5148 => "11111111",
		5149 => "11111111",
		5150 => "11110011",
		5151 => "01100100",
		5152 => "01010011",
		5153 => "11111111",
		5154 => "11111111",
		5155 => "11111111",
		5156 => "11111111",
		5157 => "11111111",
		5158 => "11111111",
		5159 => "11111111",
		5160 => "11111111",
		5161 => "11100010",
		5162 => "01011001",
		5163 => "10000001",
		5164 => "11111111",
		5165 => "11111111",
		5166 => "11111111",
		5167 => "11111111",
		5168 => "11101110",
		5169 => "10111010",
		5170 => "01011001",
		5171 => "01011110",
		5172 => "11101110",
		5173 => "11111111",
		5174 => "10000111",
		5175 => "01010011",
		5176 => "01000111",
		5177 => "01110000",
		5178 => "01011110",
		5179 => "01001101",
		5180 => "10110100",
		5181 => "11111111",
		5182 => "11111111",
		5183 => "01110101",
		5184 => "01000111",
		5185 => "01000111",
		5186 => "01100100",
		5187 => "11010111",
		5188 => "11100010",
		5189 => "10010011",
		5190 => "01000111",
		5191 => "01000111",
		5192 => "01011001",
		5193 => "01110101",
		5194 => "11010111",
		5195 => "11111001",
		5196 => "01111100",
		5197 => "01001101",
		5198 => "10010011",
		5199 => "11000000",
		5200 => "11101110",
		5201 => "11111111",
		5202 => "11111111",
		5203 => "11111111",
		5204 => "11111111",
		5205 => "01101010",
		5206 => "01011001",
		5207 => "11101110",
		5208 => "11111111",
		5209 => "11111111",
		5210 => "11111111",
		5211 => "11111111",
		5212 => "11111111",
		5213 => "11111111",
		5214 => "11111111",
		5215 => "11101110",
		5216 => "01101010",
		5217 => "01010011",
		5218 => "11011100",
		5219 => "11111111",
		5220 => "11111111",
		5221 => "11111111",
		5222 => "11111111",
		5223 => "11111111",
		5224 => "11111111",
		5225 => "11111111",
		5226 => "11111111",
		5227 => "11111111",
		5228 => "11111111",
		5229 => "11111111",
		5230 => "11111111",
		5231 => "11111111",
		5232 => "11111111",
		5233 => "11111001",
		5234 => "10111010",
		5235 => "01000111",
		5236 => "01000111",
		5237 => "01110101",
		5238 => "10101001",
		5239 => "01110000",
		5240 => "11111111",
		5241 => "11111111",
		5242 => "11111111",
		5243 => "11111111",
		5244 => "11111111",
		5245 => "11111111",
		5246 => "11111111",
		5247 => "11111111",
		5248 => "11111111",
		5249 => "11111111",
		5250 => "11111111",
		5251 => "11111111",
		5252 => "11111111",
		5253 => "11111111",
		5254 => "11111111",
		5255 => "11111111",
		5256 => "11011100",
		5257 => "01101010",
		5258 => "11101000",
		5259 => "11111111",
		5260 => "11111111",
		5261 => "11111111",
		5262 => "10111010",
		5263 => "10100011",
		5264 => "11111111",
		5265 => "11111111",
		5266 => "11111111",
		5267 => "11111111",
		5268 => "11111111",
		5269 => "11111111",
		5270 => "11111111",
		5271 => "11111111",
		5272 => "11111111",
		5273 => "11111111",
		5274 => "11111111",
		5275 => "11111111",
		5276 => "11111111",
		5277 => "11111001",
		5278 => "01101010",
		5279 => "01001101",
		5280 => "11011100",
		5281 => "11111111",
		5282 => "11111111",
		5283 => "11111111",
		5284 => "11111111",
		5285 => "11111111",
		5286 => "11111111",
		5287 => "11111111",
		5288 => "11111111",
		5289 => "11111111",
		5290 => "10101110",
		5291 => "01000111",
		5292 => "11001011",
		5293 => "11111111",
		5294 => "11111111",
		5295 => "11111111",
		5296 => "11111111",
		5297 => "11111111",
		5298 => "11100010",
		5299 => "01000111",
		5300 => "10011110",
		5301 => "01110101",
		5302 => "01011110",
		5303 => "01110101",
		5304 => "01110101",
		5305 => "01010011",
		5306 => "01000111",
		5307 => "11010001",
		5308 => "11111111",
		5309 => "11111111",
		5310 => "11111111",
		5311 => "10100011",
		5312 => "01000111",
		5313 => "01000111",
		5314 => "10011110",
		5315 => "11111111",
		5316 => "11111111",
		5317 => "11111111",
		5318 => "10101110",
		5319 => "01000111",
		5320 => "01011001",
		5321 => "01110101",
		5322 => "01000111",
		5323 => "01101010",
		5324 => "01000111",
		5325 => "11001011",
		5326 => "11111111",
		5327 => "11111111",
		5328 => "11111111",
		5329 => "11111111",
		5330 => "11111111",
		5331 => "11111111",
		5332 => "11000101",
		5333 => "01000111",
		5334 => "10101110",
		5335 => "11111111",
		5336 => "11111111",
		5337 => "11111111",
		5338 => "11111111",
		5339 => "11111111",
		5340 => "11111111",
		5341 => "11111111",
		5342 => "11111111",
		5343 => "11111111",
		5344 => "11110011",
		5345 => "01011110",
		5346 => "01011001",
		5347 => "11101110",
		5348 => "11111111",
		5349 => "11111111",
		5350 => "11111111",
		5351 => "11111111",
		5352 => "11111111",
		5353 => "11111111",
		5354 => "11111111",
		5355 => "11111001",
		5356 => "11111001",
		5357 => "11111111",
		5358 => "11111111",
		5359 => "11101110",
		5360 => "10100011",
		5361 => "01011001",
		5362 => "01000111",
		5363 => "10000111",
		5364 => "11010111",
		5365 => "11111111",
		5366 => "11111111",
		5367 => "11010111",
		5368 => "11111001",
		5369 => "11111111",
		5370 => "11111111",
		5371 => "11111111",
		5372 => "11111111",
		5373 => "11111111",
		5374 => "11111111",
		5375 => "11111111",
		5376 => "11111111",
		5377 => "11111111",
		5378 => "11111111",
		5379 => "11111111",
		5380 => "11111111",
		5381 => "11111111",
		5382 => "11111111",
		5383 => "11111111",
		5384 => "10000001",
		5385 => "01000111",
		5386 => "01000111",
		5387 => "01111100",
		5388 => "11001011",
		5389 => "11111111",
		5390 => "10001100",
		5391 => "11010001",
		5392 => "11111111",
		5393 => "11111111",
		5394 => "11111111",
		5395 => "11111111",
		5396 => "11111111",
		5397 => "11111111",
		5398 => "11111111",
		5399 => "11111111",
		5400 => "11111111",
		5401 => "11111111",
		5402 => "11111111",
		5403 => "11111111",
		5404 => "11111111",
		5405 => "10100011",
		5406 => "01000111",
		5407 => "11001011",
		5408 => "11111111",
		5409 => "11111111",
		5410 => "11111111",
		5411 => "11111111",
		5412 => "11111111",
		5413 => "11111111",
		5414 => "11111111",
		5415 => "11111111",
		5416 => "11111111",
		5417 => "11111111",
		5418 => "11111001",
		5419 => "01100100",
		5420 => "01111100",
		5421 => "11111111",
		5422 => "11111111",
		5423 => "11111111",
		5424 => "11111111",
		5425 => "11111111",
		5426 => "11111111",
		5427 => "01000111",
		5428 => "01000111",
		5429 => "01001101",
		5430 => "11111111",
		5431 => "11111111",
		5432 => "11110011",
		5433 => "01001101",
		5434 => "10000001",
		5435 => "11111111",
		5436 => "11111111",
		5437 => "11111111",
		5438 => "11101110",
		5439 => "01100100",
		5440 => "01000111",
		5441 => "01000111",
		5442 => "01101010",
		5443 => "11111111",
		5444 => "11111111",
		5445 => "11111111",
		5446 => "11111111",
		5447 => "01111100",
		5448 => "01011001",
		5449 => "11111001",
		5450 => "10000111",
		5451 => "01000111",
		5452 => "01010011",
		5453 => "11111111",
		5454 => "11111111",
		5455 => "11111111",
		5456 => "11111111",
		5457 => "11111111",
		5458 => "11111111",
		5459 => "11111111",
		5460 => "01111100",
		5461 => "01011110",
		5462 => "11111111",
		5463 => "11111111",
		5464 => "11111111",
		5465 => "11111111",
		5466 => "11111111",
		5467 => "11111111",
		5468 => "11111111",
		5469 => "11111111",
		5470 => "11111111",
		5471 => "11111111",
		5472 => "11111111",
		5473 => "11101000",
		5474 => "01010011",
		5475 => "10000111",
		5476 => "11111111",
		5477 => "11111111",
		5478 => "11111111",
		5479 => "11111111",
		5480 => "11111111",
		5481 => "11111111",
		5482 => "11111111",
		5483 => "11011100",
		5484 => "01110101",
		5485 => "11011100",
		5486 => "10001100",
		5487 => "01001101",
		5488 => "01000111",
		5489 => "01010011",
		5490 => "10011000",
		5491 => "11111111",
		5492 => "11111111",
		5493 => "11111111",
		5494 => "11111111",
		5495 => "11111111",
		5496 => "11111111",
		5497 => "11111111",
		5498 => "11111111",
		5499 => "11111111",
		5500 => "11111111",
		5501 => "11111111",
		5502 => "11111111",
		5503 => "11111111",
		5504 => "11111111",
		5505 => "11111111",
		5506 => "11111111",
		5507 => "11111111",
		5508 => "11111111",
		5509 => "11111111",
		5510 => "11111111",
		5511 => "11101110",
		5512 => "01100100",
		5513 => "10110100",
		5514 => "01110000",
		5515 => "01000111",
		5516 => "01000111",
		5517 => "10110100",
		5518 => "01110101",
		5519 => "11111111",
		5520 => "11111111",
		5521 => "11111111",
		5522 => "11111111",
		5523 => "11111111",
		5524 => "11111111",
		5525 => "11111111",
		5526 => "11111111",
		5527 => "11111111",
		5528 => "11111111",
		5529 => "11111111",
		5530 => "11111111",
		5531 => "11111111",
		5532 => "11011100",
		5533 => "01001101",
		5534 => "10010011",
		5535 => "11111111",
		5536 => "11111111",
		5537 => "11111111",
		5538 => "11111111",
		5539 => "11111111",
		5540 => "11111111",
		5541 => "11111111",
		5542 => "11111111",
		5543 => "11111111",
		5544 => "11111111",
		5545 => "11111111",
		5546 => "11111111",
		5547 => "10011110",
		5548 => "01001101",
		5549 => "11110011",
		5550 => "11111111",
		5551 => "11111111",
		5552 => "11111111",
		5553 => "11111111",
		5554 => "11011100",
		5555 => "01000111",
		5556 => "01000111",
		5557 => "10111010",
		5558 => "11111111",
		5559 => "11111111",
		5560 => "11001011",
		5561 => "01000111",
		5562 => "11000101",
		5563 => "11111111",
		5564 => "11111111",
		5565 => "10100011",
		5566 => "01001101",
		5567 => "01000111",
		5568 => "10011000",
		5569 => "01000111",
		5570 => "01000111",
		5571 => "01101010",
		5572 => "11010111",
		5573 => "11111111",
		5574 => "11111111",
		5575 => "11010001",
		5576 => "01000111",
		5577 => "11000101",
		5578 => "11111001",
		5579 => "01100100",
		5580 => "01000111",
		5581 => "11101000",
		5582 => "11111111",
		5583 => "11111111",
		5584 => "11111111",
		5585 => "11111111",
		5586 => "11111111",
		5587 => "11110011",
		5588 => "01001101",
		5589 => "10011110",
		5590 => "11111111",
		5591 => "11111111",
		5592 => "11111111",
		5593 => "11111111",
		5594 => "11111111",
		5595 => "11111111",
		5596 => "11111111",
		5597 => "11111111",
		5598 => "11111111",
		5599 => "11111111",
		5600 => "11111111",
		5601 => "11111111",
		5602 => "10111010",
		5603 => "01000111",
		5604 => "11000000",
		5605 => "11111111",
		5606 => "11111111",
		5607 => "11111111",
		5608 => "11111111",
		5609 => "11111111",
		5610 => "11111111",
		5611 => "11111111",
		5612 => "10000001",
		5613 => "01000111",
		5614 => "01000111",
		5615 => "01011001",
		5616 => "10101001",
		5617 => "11110011",
		5618 => "11111111",
		5619 => "11111111",
		5620 => "11111111",
		5621 => "11111111",
		5622 => "11111111",
		5623 => "11111111",
		5624 => "11111111",
		5625 => "11111111",
		5626 => "11111111",
		5627 => "11111111",
		5628 => "11111111",
		5629 => "11111111",
		5630 => "11111111",
		5631 => "11111111",
		5632 => "11111111",
		5633 => "11111111",
		5634 => "11111111",
		5635 => "11111111",
		5636 => "11111111",
		5637 => "11111111",
		5638 => "11111111",
		5639 => "11101000",
		5640 => "11101000",
		5641 => "11111111",
		5642 => "11111111",
		5643 => "11010111",
		5644 => "10001100",
		5645 => "01000111",
		5646 => "01010011",
		5647 => "10010011",
		5648 => "11101000",
		5649 => "11111111",
		5650 => "11111111",
		5651 => "10111010",
		5652 => "11100010",
		5653 => "11111111",
		5654 => "11111111",
		5655 => "11111111",
		5656 => "11111111",
		5657 => "11111111",
		5658 => "11111111",
		5659 => "11111111",
		5660 => "01101010",
		5661 => "01011110",
		5662 => "11111001",
		5663 => "11111111",
		5664 => "11111111",
		5665 => "11111111",
		5666 => "11111111",
		5667 => "11111111",
		5668 => "11111111",
		5669 => "11111111",
		5670 => "11111111",
		5671 => "11111111",
		5672 => "11111111",
		5673 => "11111111",
		5674 => "11111111",
		5675 => "11000101",
		5676 => "01000111",
		5677 => "11010001",
		5678 => "11111111",
		5679 => "11111111",
		5680 => "11111111",
		5681 => "11111111",
		5682 => "10011000",
		5683 => "01000111",
		5684 => "01100100",
		5685 => "11111111",
		5686 => "11100010",
		5687 => "11101110",
		5688 => "10110100",
		5689 => "01000111",
		5690 => "11101110",
		5691 => "11111111",
		5692 => "10101001",
		5693 => "01000111",
		5694 => "01011110",
		5695 => "01000111",
		5696 => "11010111",
		5697 => "01000111",
		5698 => "01011001",
		5699 => "01011110",
		5700 => "01001101",
		5701 => "11001011",
		5702 => "11111111",
		5703 => "11101110",
		5704 => "01000111",
		5705 => "10101110",
		5706 => "11111111",
		5707 => "11001011",
		5708 => "01000111",
		5709 => "01110101",
		5710 => "11101110",
		5711 => "11111111",
		5712 => "11111111",
		5713 => "11111111",
		5714 => "11111111",
		5715 => "11010111",
		5716 => "01000111",
		5717 => "11000101",
		5718 => "11111111",
		5719 => "11111111",
		5720 => "11111111",
		5721 => "11111111",
		5722 => "11111111",
		5723 => "11111111",
		5724 => "11111111",
		5725 => "11111111",
		5726 => "11111111",
		5727 => "11111111",
		5728 => "11111111",
		5729 => "11111111",
		5730 => "11111111",
		5731 => "01111100",
		5732 => "01011001",
		5733 => "11111001",
		5734 => "11111111",
		5735 => "11111111",
		5736 => "11111111",
		5737 => "11111111",
		5738 => "11111111",
		5739 => "11111111",
		5740 => "11011100",
		5741 => "01000111",
		5742 => "10101110",
		5743 => "11111111",
		5744 => "11111111",
		5745 => "11111111",
		5746 => "11111111",
		5747 => "11111111",
		5748 => "11111111",
		5749 => "11111111",
		5750 => "11111111",
		5751 => "11010001",
		5752 => "10100011",
		5753 => "10100011",
		5754 => "11111111",
		5755 => "11111111",
		5756 => "11111111",
		5757 => "11111111",
		5758 => "11111111",
		5759 => "11111111",
		5760 => "11111111",
		5761 => "11111111",
		5762 => "11111111",
		5763 => "11111111",
		5764 => "11111111",
		5765 => "11111111",
		5766 => "11111111",
		5767 => "11111111",
		5768 => "11111111",
		5769 => "11111111",
		5770 => "11111111",
		5771 => "11111111",
		5772 => "11111111",
		5773 => "10100011",
		5774 => "01011001",
		5775 => "01000111",
		5776 => "01000111",
		5777 => "01111100",
		5778 => "10011110",
		5779 => "01101010",
		5780 => "11111111",
		5781 => "11111111",
		5782 => "11111111",
		5783 => "11111111",
		5784 => "11111111",
		5785 => "11111111",
		5786 => "11111111",
		5787 => "11010001",
		5788 => "01000111",
		5789 => "10001100",
		5790 => "11111111",
		5791 => "11111111",
		5792 => "11111111",
		5793 => "11111111",
		5794 => "11111111",
		5795 => "11111111",
		5796 => "11111111",
		5797 => "11111111",
		5798 => "11111111",
		5799 => "11111111",
		5800 => "11111111",
		5801 => "11111111",
		5802 => "11111111",
		5803 => "11101110",
		5804 => "01000111",
		5805 => "10100011",
		5806 => "11111111",
		5807 => "11111111",
		5808 => "11111111",
		5809 => "10101001",
		5810 => "01000111",
		5811 => "01000111",
		5812 => "10001100",
		5813 => "11111111",
		5814 => "01000111",
		5815 => "10001100",
		5816 => "10011000",
		5817 => "01010011",
		5818 => "11111111",
		5819 => "11111111",
		5820 => "01010011",
		5821 => "01010011",
		5822 => "10011110",
		5823 => "01000111",
		5824 => "10001100",
		5825 => "11001011",
		5826 => "11101110",
		5827 => "11001011",
		5828 => "01000111",
		5829 => "01100100",
		5830 => "11111111",
		5831 => "11111111",
		5832 => "01011001",
		5833 => "10010011",
		5834 => "01011110",
		5835 => "11000101",
		5836 => "01000111",
		5837 => "01000111",
		5838 => "01010011",
		5839 => "11101110",
		5840 => "11111111",
		5841 => "11111111",
		5842 => "11111111",
		5843 => "10101001",
		5844 => "01000111",
		5845 => "11101000",
		5846 => "11111111",
		5847 => "11111111",
		5848 => "11111111",
		5849 => "11111111",
		5850 => "11111111",
		5851 => "11111111",
		5852 => "11111111",
		5853 => "11111111",
		5854 => "11111111",
		5855 => "11111111",
		5856 => "11111111",
		5857 => "11111111",
		5858 => "11111111",
		5859 => "10011110",
		5860 => "01000111",
		5861 => "10110100",
		5862 => "11111111",
		5863 => "11111111",
		5864 => "11111111",
		5865 => "11111111",
		5866 => "11111111",
		5867 => "11111111",
		5868 => "11111111",
		5869 => "01110101",
		5870 => "11101000",
		5871 => "11111111",
		5872 => "11111111",
		5873 => "11111111",
		5874 => "11111111",
		5875 => "11111111",
		5876 => "11111111",
		5877 => "11111111",
		5878 => "11000101",
		5879 => "01110101",
		5880 => "01011110",
		5881 => "01011001",
		5882 => "11111111",
		5883 => "11111111",
		5884 => "11111111",
		5885 => "11111111",
		5886 => "11111111",
		5887 => "11111111",
		5888 => "11111111",
		5889 => "11111111",
		5890 => "11111111",
		5891 => "11111111",
		5892 => "11111111",
		5893 => "11111111",
		5894 => "11111111",
		5895 => "11111111",
		5896 => "11111111",
		5897 => "11111111",
		5898 => "11111111",
		5899 => "11111111",
		5900 => "11111111",
		5901 => "11111111",
		5902 => "11111111",
		5903 => "10111010",
		5904 => "01110000",
		5905 => "01000111",
		5906 => "01000111",
		5907 => "10111010",
		5908 => "11111111",
		5909 => "11111111",
		5910 => "11111111",
		5911 => "11111111",
		5912 => "11111111",
		5913 => "11111111",
		5914 => "11111111",
		5915 => "10000001",
		5916 => "01000111",
		5917 => "01011001",
		5918 => "11111111",
		5919 => "11111111",
		5920 => "11111111",
		5921 => "11111111",
		5922 => "11111111",
		5923 => "11111111",
		5924 => "11111111",
		5925 => "11111111",
		5926 => "11111111",
		5927 => "11111111",
		5928 => "11111111",
		5929 => "11111111",
		5930 => "11111111",
		5931 => "11111111",
		5932 => "01101010",
		5933 => "01011001",
		5934 => "11111111",
		5935 => "11111111",
		5936 => "11101110",
		5937 => "01001101",
		5938 => "01111100",
		5939 => "01011110",
		5940 => "10001100",
		5941 => "11000101",
		5942 => "01000111",
		5943 => "01100100",
		5944 => "01100100",
		5945 => "01110000",
		5946 => "11111111",
		5947 => "11011100",
		5948 => "01000111",
		5949 => "01000111",
		5950 => "01000111",
		5951 => "01000111",
		5952 => "01000111",
		5953 => "01101010",
		5954 => "10100011",
		5955 => "01110000",
		5956 => "01000111",
		5957 => "01000111",
		5958 => "11011100",
		5959 => "11111111",
		5960 => "01111100",
		5961 => "01100100",
		5962 => "01000111",
		5963 => "01000111",
		5964 => "01000111",
		5965 => "10000111",
		5966 => "01001101",
		5967 => "10011000",
		5968 => "11111111",
		5969 => "11111111",
		5970 => "11111111",
		5971 => "01100100",
		5972 => "01101010",
		5973 => "11111111",
		5974 => "11111111",
		5975 => "11111111",
		5976 => "11111111",
		5977 => "11111111",
		5978 => "11111111",
		5979 => "11111111",
		5980 => "11111111",
		5981 => "11111111",
		5982 => "11111111",
		5983 => "11111111",
		5984 => "11111111",
		5985 => "11111111",
		5986 => "11111111",
		5987 => "01111100",
		5988 => "01000111",
		5989 => "01101010",
		5990 => "11111111",
		5991 => "11111111",
		5992 => "11111111",
		5993 => "11111111",
		5994 => "11111111",
		5995 => "11111111",
		5996 => "11111111",
		5997 => "11011100",
		5998 => "11111001",
		5999 => "11111111",
		6000 => "11111111",
		6001 => "11111111",
		6002 => "11111111",
		6003 => "11111111",
		6004 => "11111111",
		6005 => "11111111",
		6006 => "11111111",
		6007 => "11111111",
		6008 => "11111111",
		6009 => "01111100",
		6010 => "11011100",
		6011 => "11111111",
		6012 => "11111111",
		6013 => "11111111",
		6014 => "11111111",
		6015 => "11111111",
		6016 => "11111111",
		6017 => "11111111",
		6018 => "11111111",
		6019 => "11111111",
		6020 => "11111111",
		6021 => "11111111",
		6022 => "11111111",
		6023 => "11111111",
		6024 => "11111111",
		6025 => "11111111",
		6026 => "11111111",
		6027 => "11111111",
		6028 => "11111111",
		6029 => "11111111",
		6030 => "11111111",
		6031 => "11111111",
		6032 => "11111111",
		6033 => "10111010",
		6034 => "01011001",
		6035 => "11111001",
		6036 => "11111111",
		6037 => "11111111",
		6038 => "11111111",
		6039 => "11111111",
		6040 => "11111111",
		6041 => "11111111",
		6042 => "11101000",
		6043 => "01000111",
		6044 => "01101010",
		6045 => "01000111",
		6046 => "10110100",
		6047 => "11111111",
		6048 => "11111111",
		6049 => "11111111",
		6050 => "11111111",
		6051 => "11111111",
		6052 => "11111111",
		6053 => "11111111",
		6054 => "11111111",
		6055 => "11111111",
		6056 => "11111111",
		6057 => "11111111",
		6058 => "11111111",
		6059 => "11111111",
		6060 => "11000101",
		6061 => "01000111",
		6062 => "10101110",
		6063 => "11111111",
		6064 => "10101110",
		6065 => "01000111",
		6066 => "11011100",
		6067 => "01010011",
		6068 => "10100011",
		6069 => "10011110",
		6070 => "10111010",
		6071 => "01000111",
		6072 => "01000111",
		6073 => "11010111",
		6074 => "11111111",
		6075 => "10111010",
		6076 => "01000111",
		6077 => "11011100",
		6078 => "11001011",
		6079 => "11000000",
		6080 => "01011001",
		6081 => "01000111",
		6082 => "01000111",
		6083 => "01000111",
		6084 => "01000111",
		6085 => "01000111",
		6086 => "10111010",
		6087 => "11111111",
		6088 => "11001011",
		6089 => "01000111",
		6090 => "10000001",
		6091 => "01000111",
		6092 => "01000111",
		6093 => "10011110",
		6094 => "10010011",
		6095 => "01001101",
		6096 => "11111001",
		6097 => "11111111",
		6098 => "10101001",
		6099 => "01000111",
		6100 => "11000101",
		6101 => "11111111",
		6102 => "11111111",
		6103 => "11111111",
		6104 => "11111111",
		6105 => "11111111",
		6106 => "11111111",
		6107 => "11111111",
		6108 => "11111111",
		6109 => "11111111",
		6110 => "11101110",
		6111 => "11100010",
		6112 => "11111111",
		6113 => "11111001",
		6114 => "10101001",
		6115 => "01000111",
		6116 => "10000001",
		6117 => "01000111",
		6118 => "11001011",
		6119 => "11111111",
		6120 => "11111111",
		6121 => "11111111",
		6122 => "11111111",
		6123 => "11111111",
		6124 => "11111111",
		6125 => "11111111",
		6126 => "11111111",
		6127 => "11111111",
		6128 => "11111111",
		6129 => "11111111",
		6130 => "11111111",
		6131 => "11111111",
		6132 => "11111111",
		6133 => "11111111",
		6134 => "11111111",
		6135 => "11111111",
		6136 => "11111111",
		6137 => "10101110",
		6138 => "10101001",
		6139 => "11111111",
		6140 => "11111111",
		6141 => "11111111",
		6142 => "11111111",
		6143 => "11111111",
		6144 => "11111111",
		6145 => "11111111",
		6146 => "11111111",
		6147 => "11111111",
		6148 => "11111111",
		6149 => "11111111",
		6150 => "10010011",
		6151 => "11111111",
		6152 => "11111111",
		6153 => "11111111",
		6154 => "11111111",
		6155 => "11111111",
		6156 => "11111111",
		6157 => "11111111",
		6158 => "11111111",
		6159 => "11111111",
		6160 => "11111111",
		6161 => "11010001",
		6162 => "10101001",
		6163 => "11111111",
		6164 => "11111111",
		6165 => "11111111",
		6166 => "11111111",
		6167 => "11111111",
		6168 => "11111111",
		6169 => "11111111",
		6170 => "10011000",
		6171 => "01001101",
		6172 => "11110011",
		6173 => "01110101",
		6174 => "01000111",
		6175 => "01011110",
		6176 => "10000111",
		6177 => "10011110",
		6178 => "11111111",
		6179 => "11111111",
		6180 => "11111111",
		6181 => "11111111",
		6182 => "11111111",
		6183 => "11111111",
		6184 => "11111111",
		6185 => "11111111",
		6186 => "11111111",
		6187 => "11111111",
		6188 => "11111111",
		6189 => "10000001",
		6190 => "01001101",
		6191 => "11011100",
		6192 => "10000111",
		6193 => "01010011",
		6194 => "10110100",
		6195 => "01000111",
		6196 => "10111010",
		6197 => "10101001",
		6198 => "11110011",
		6199 => "11101000",
		6200 => "11111001",
		6201 => "11111111",
		6202 => "11111111",
		6203 => "10000001",
		6204 => "01000111",
		6205 => "11101000",
		6206 => "11111111",
		6207 => "10111010",
		6208 => "01000111",
		6209 => "10000001",
		6210 => "01110000",
		6211 => "01000111",
		6212 => "10001100",
		6213 => "01001101",
		6214 => "10010011",
		6215 => "11111111",
		6216 => "11111111",
		6217 => "11001011",
		6218 => "11111001",
		6219 => "01011001",
		6220 => "01000111",
		6221 => "01110101",
		6222 => "01110000",
		6223 => "01000111",
		6224 => "11011100",
		6225 => "11000101",
		6226 => "01000111",
		6227 => "10000111",
		6228 => "11111111",
		6229 => "11111111",
		6230 => "11111111",
		6231 => "11111111",
		6232 => "11111111",
		6233 => "11111111",
		6234 => "11111111",
		6235 => "11111111",
		6236 => "11111111",
		6237 => "11111111",
		6238 => "10000001",
		6239 => "01000111",
		6240 => "01110000",
		6241 => "01010011",
		6242 => "01000111",
		6243 => "10000111",
		6244 => "11111111",
		6245 => "01011001",
		6246 => "10000001",
		6247 => "11111111",
		6248 => "11111111",
		6249 => "11111111",
		6250 => "11111111",
		6251 => "11111111",
		6252 => "11111111",
		6253 => "11111111",
		6254 => "11111111",
		6255 => "11111111",
		6256 => "11111111",
		6257 => "11111111",
		6258 => "11111111",
		6259 => "11111111",
		6260 => "11111111",
		6261 => "11111111",
		6262 => "11111111",
		6263 => "11111111",
		6264 => "11111001",
		6265 => "10110100",
		6266 => "01110101",
		6267 => "11111111",
		6268 => "11111111",
		6269 => "11111111",
		6270 => "11111111",
		6271 => "11111111",
		6272 => "11111111",
		6273 => "11111111",
		6274 => "11111111",
		6275 => "11111111",
		6276 => "11111111",
		6277 => "11101110",
		6278 => "01010011",
		6279 => "11100010",
		6280 => "11111111",
		6281 => "11111111",
		6282 => "11111111",
		6283 => "11111111",
		6284 => "11111111",
		6285 => "11111111",
		6286 => "11111111",
		6287 => "11111111",
		6288 => "11111111",
		6289 => "11111111",
		6290 => "11110011",
		6291 => "11111111",
		6292 => "11111111",
		6293 => "11111111",
		6294 => "11111111",
		6295 => "11111111",
		6296 => "11111111",
		6297 => "11111111",
		6298 => "01010011",
		6299 => "10000001",
		6300 => "11111111",
		6301 => "11110011",
		6302 => "10011110",
		6303 => "01101010",
		6304 => "01011001",
		6305 => "01001101",
		6306 => "11101110",
		6307 => "11111111",
		6308 => "11111111",
		6309 => "11101000",
		6310 => "10010011",
		6311 => "11101000",
		6312 => "11111111",
		6313 => "11111111",
		6314 => "11111111",
		6315 => "11111111",
		6316 => "11111111",
		6317 => "11110011",
		6318 => "01011001",
		6319 => "01010011",
		6320 => "01011110",
		6321 => "01000111",
		6322 => "01000111",
		6323 => "01000111",
		6324 => "11011100",
		6325 => "10000111",
		6326 => "10100011",
		6327 => "11111111",
		6328 => "11111111",
		6329 => "11111111",
		6330 => "11000101",
		6331 => "01000111",
		6332 => "01000111",
		6333 => "01011001",
		6334 => "01110101",
		6335 => "01000111",
		6336 => "01000111",
		6337 => "01001101",
		6338 => "11101110",
		6339 => "11101000",
		6340 => "11111111",
		6341 => "01101010",
		6342 => "01001101",
		6343 => "11101000",
		6344 => "11111111",
		6345 => "11111111",
		6346 => "11011100",
		6347 => "01000111",
		6348 => "01010011",
		6349 => "01000111",
		6350 => "01000111",
		6351 => "01000111",
		6352 => "10001100",
		6353 => "01001101",
		6354 => "01110000",
		6355 => "11111001",
		6356 => "11111111",
		6357 => "11111111",
		6358 => "11111111",
		6359 => "11111111",
		6360 => "11111111",
		6361 => "11101000",
		6362 => "01110000",
		6363 => "11010001",
		6364 => "11111111",
		6365 => "11111111",
		6366 => "01000111",
		6367 => "10000001",
		6368 => "01110101",
		6369 => "01110101",
		6370 => "10101110",
		6371 => "11111111",
		6372 => "11111111",
		6373 => "10010011",
		6374 => "01000111",
		6375 => "11110011",
		6376 => "11111111",
		6377 => "11111111",
		6378 => "11111111",
		6379 => "11111111",
		6380 => "11111111",
		6381 => "11111111",
		6382 => "11111111",
		6383 => "11100010",
		6384 => "11111111",
		6385 => "11111111",
		6386 => "11111111",
		6387 => "11111111",
		6388 => "11111111",
		6389 => "11010111",
		6390 => "10101001",
		6391 => "01110101",
		6392 => "01000111",
		6393 => "01000111",
		6394 => "01001101",
		6395 => "11111001",
		6396 => "11111111",
		6397 => "11111111",
		6398 => "11111111",
		6399 => "11111111",
		6400 => "11111111",
		6401 => "11111111",
		6402 => "11111111",
		6403 => "11111111",
		6404 => "11111111",
		6405 => "11001011",
		6406 => "01000111",
		6407 => "01000111",
		6408 => "01000111",
		6409 => "01110101",
		6410 => "10011000",
		6411 => "10111010",
		6412 => "11010111",
		6413 => "11111111",
		6414 => "11111111",
		6415 => "11111111",
		6416 => "11111111",
		6417 => "11111111",
		6418 => "11111111",
		6419 => "11111111",
		6420 => "11111111",
		6421 => "11111111",
		6422 => "11111111",
		6423 => "11111111",
		6424 => "11111111",
		6425 => "11011100",
		6426 => "01000111",
		6427 => "11000000",
		6428 => "11111111",
		6429 => "11111111",
		6430 => "11111111",
		6431 => "11111111",
		6432 => "11111111",
		6433 => "01010011",
		6434 => "01101010",
		6435 => "10110100",
		6436 => "10101001",
		6437 => "01011001",
		6438 => "01000111",
		6439 => "10101001",
		6440 => "11111111",
		6441 => "11111111",
		6442 => "11111111",
		6443 => "11111111",
		6444 => "11111111",
		6445 => "11011100",
		6446 => "01000111",
		6447 => "01000111",
		6448 => "01000111",
		6449 => "10011110",
		6450 => "10000001",
		6451 => "10111010",
		6452 => "10101110",
		6453 => "01000111",
		6454 => "01000111",
		6455 => "01110000",
		6456 => "10100011",
		6457 => "10000001",
		6458 => "01000111",
		6459 => "01000111",
		6460 => "01100100",
		6461 => "01000111",
		6462 => "01000111",
		6463 => "01111100",
		6464 => "11010001",
		6465 => "01001101",
		6466 => "01011110",
		6467 => "10110100",
		6468 => "10010011",
		6469 => "01000111",
		6470 => "01000111",
		6471 => "01011001",
		6472 => "10101001",
		6473 => "11010001",
		6474 => "01011001",
		6475 => "01000111",
		6476 => "01101010",
		6477 => "10000001",
		6478 => "10011110",
		6479 => "01100100",
		6480 => "01000111",
		6481 => "01000111",
		6482 => "01110000",
		6483 => "11111111",
		6484 => "11111111",
		6485 => "11111111",
		6486 => "11111111",
		6487 => "11111111",
		6488 => "11111111",
		6489 => "10101110",
		6490 => "01000111",
		6491 => "01001101",
		6492 => "10001100",
		6493 => "10010011",
		6494 => "01100100",
		6495 => "11111001",
		6496 => "11111111",
		6497 => "11111111",
		6498 => "11111111",
		6499 => "11111111",
		6500 => "11111111",
		6501 => "11010001",
		6502 => "01000111",
		6503 => "11000101",
		6504 => "11111111",
		6505 => "11111111",
		6506 => "11111111",
		6507 => "11111111",
		6508 => "11111111",
		6509 => "11111111",
		6510 => "11111111",
		6511 => "01110000",
		6512 => "11101110",
		6513 => "11111111",
		6514 => "11100010",
		6515 => "10000001",
		6516 => "01010011",
		6517 => "01000111",
		6518 => "01000111",
		6519 => "01000111",
		6520 => "01101010",
		6521 => "10011110",
		6522 => "01111100",
		6523 => "11000101",
		6524 => "11111111",
		6525 => "11111111",
		6526 => "11111111",
		6527 => "11111111",
		6528 => "11111111",
		6529 => "11111111",
		6530 => "11111111",
		6531 => "11111111",
		6532 => "11111111",
		6533 => "10101001",
		6534 => "10110100",
		6535 => "11100010",
		6536 => "11000101",
		6537 => "10100011",
		6538 => "01111100",
		6539 => "01011110",
		6540 => "01000111",
		6541 => "01110101",
		6542 => "10111010",
		6543 => "11110011",
		6544 => "11111111",
		6545 => "11111111",
		6546 => "11111111",
		6547 => "11111111",
		6548 => "11111111",
		6549 => "11111111",
		6550 => "11111111",
		6551 => "11111111",
		6552 => "11111111",
		6553 => "10101110",
		6554 => "01001101",
		6555 => "11111001",
		6556 => "11111111",
		6557 => "11111111",
		6558 => "11111111",
		6559 => "11111111",
		6560 => "11111111",
		6561 => "11000101",
		6562 => "01101010",
		6563 => "01000111",
		6564 => "01010011",
		6565 => "10001100",
		6566 => "01101010",
		6567 => "01101010",
		6568 => "11111111",
		6569 => "11111111",
		6570 => "11111111",
		6571 => "11010001",
		6572 => "01110101",
		6573 => "10100011",
		6574 => "01000111",
		6575 => "01000111",
		6576 => "01000111",
		6577 => "11100010",
		6578 => "11111111",
		6579 => "11111111",
		6580 => "01100100",
		6581 => "01000111",
		6582 => "01110000",
		6583 => "01010011",
		6584 => "01000111",
		6585 => "01011110",
		6586 => "10101001",
		6587 => "10011110",
		6588 => "01000111",
		6589 => "01011001",
		6590 => "10001100",
		6591 => "11111001",
		6592 => "11111111",
		6593 => "11010001",
		6594 => "01101010",
		6595 => "01000111",
		6596 => "01000111",
		6597 => "10011110",
		6598 => "11100010",
		6599 => "01110000",
		6600 => "01000111",
		6601 => "01000111",
		6602 => "01100100",
		6603 => "10000001",
		6604 => "01001101",
		6605 => "11111001",
		6606 => "11111111",
		6607 => "10011000",
		6608 => "01000111",
		6609 => "01000111",
		6610 => "01000111",
		6611 => "11110011",
		6612 => "01001101",
		6613 => "10111010",
		6614 => "11111111",
		6615 => "11111111",
		6616 => "11110011",
		6617 => "01011110",
		6618 => "01110000",
		6619 => "10001100",
		6620 => "01000111",
		6621 => "01010011",
		6622 => "11011100",
		6623 => "11111111",
		6624 => "11111111",
		6625 => "11111111",
		6626 => "11111111",
		6627 => "11111111",
		6628 => "11111111",
		6629 => "11111111",
		6630 => "01010011",
		6631 => "10010011",
		6632 => "11111111",
		6633 => "11111111",
		6634 => "11111111",
		6635 => "11111111",
		6636 => "11111111",
		6637 => "11111111",
		6638 => "11111111",
		6639 => "10010011",
		6640 => "01100100",
		6641 => "01011110",
		6642 => "01000111",
		6643 => "01000111",
		6644 => "01011110",
		6645 => "10010011",
		6646 => "11000000",
		6647 => "11110011",
		6648 => "11111111",
		6649 => "11111111",
		6650 => "10111010",
		6651 => "10011000",
		6652 => "11111111",
		6653 => "11111111",
		6654 => "11111111",
		6655 => "11111111",
		6656 => "11111111",
		6657 => "11111111",
		6658 => "11111111",
		6659 => "11111111",
		6660 => "11111111",
		6661 => "11100010",
		6662 => "11111111",
		6663 => "11111111",
		6664 => "11111111",
		6665 => "11111111",
		6666 => "11111111",
		6667 => "11111111",
		6668 => "11111001",
		6669 => "10101110",
		6670 => "01110000",
		6671 => "01110000",
		6672 => "11111001",
		6673 => "11111111",
		6674 => "11111111",
		6675 => "11111111",
		6676 => "11111111",
		6677 => "11111111",
		6678 => "11111111",
		6679 => "11111111",
		6680 => "11111111",
		6681 => "01111100",
		6682 => "01000111",
		6683 => "11010001",
		6684 => "11111111",
		6685 => "11111111",
		6686 => "11111111",
		6687 => "11111111",
		6688 => "11111111",
		6689 => "11111111",
		6690 => "11111111",
		6691 => "11101110",
		6692 => "11111111",
		6693 => "11111111",
		6694 => "11101000",
		6695 => "01010011",
		6696 => "01110000",
		6697 => "10100011",
		6698 => "10011000",
		6699 => "01001101",
		6700 => "01101010",
		6701 => "11010111",
		6702 => "01000111",
		6703 => "01100100",
		6704 => "01000111",
		6705 => "10101110",
		6706 => "11111111",
		6707 => "11100010",
		6708 => "01000111",
		6709 => "01000111",
		6710 => "01011001",
		6711 => "01000111",
		6712 => "11000101",
		6713 => "11111111",
		6714 => "11111111",
		6715 => "11111111",
		6716 => "11111111",
		6717 => "11111111",
		6718 => "11111111",
		6719 => "11111111",
		6720 => "11111111",
		6721 => "11111111",
		6722 => "11111111",
		6723 => "11101000",
		6724 => "11111111",
		6725 => "11111111",
		6726 => "11111111",
		6727 => "11111111",
		6728 => "01111100",
		6729 => "01000111",
		6730 => "10010011",
		6731 => "10100011",
		6732 => "01000111",
		6733 => "11101110",
		6734 => "11111111",
		6735 => "10011110",
		6736 => "01000111",
		6737 => "01100100",
		6738 => "01101010",
		6739 => "11111001",
		6740 => "10001100",
		6741 => "01000111",
		6742 => "01111100",
		6743 => "10011110",
		6744 => "01011110",
		6745 => "01011001",
		6746 => "11101000",
		6747 => "11111111",
		6748 => "11111111",
		6749 => "11111111",
		6750 => "11111111",
		6751 => "11111111",
		6752 => "11111111",
		6753 => "11111111",
		6754 => "11111111",
		6755 => "11111111",
		6756 => "11111111",
		6757 => "11101110",
		6758 => "01001101",
		6759 => "01011110",
		6760 => "11111111",
		6761 => "11111111",
		6762 => "11111111",
		6763 => "11111111",
		6764 => "11111111",
		6765 => "11111111",
		6766 => "11111111",
		6767 => "11000101",
		6768 => "01000111",
		6769 => "01010011",
		6770 => "10000001",
		6771 => "11101000",
		6772 => "11111111",
		6773 => "11111111",
		6774 => "11111111",
		6775 => "11111111",
		6776 => "11111111",
		6777 => "11111111",
		6778 => "11110011",
		6779 => "01100100",
		6780 => "11111111",
		6781 => "11111111",
		6782 => "11111111",
		6783 => "11111111",
		6784 => "11111111",
		6785 => "11111111",
		6786 => "11111111",
		6787 => "11111111",
		6788 => "11111111",
		6789 => "11111111",
		6790 => "11111111",
		6791 => "11111111",
		6792 => "11111111",
		6793 => "11111111",
		6794 => "11111111",
		6795 => "11111111",
		6796 => "11111111",
		6797 => "11111111",
		6798 => "11111111",
		6799 => "10010011",
		6800 => "10011110",
		6801 => "11111111",
		6802 => "11111111",
		6803 => "11111111",
		6804 => "11111111",
		6805 => "11111111",
		6806 => "11111111",
		6807 => "11111111",
		6808 => "11111001",
		6809 => "01001101",
		6810 => "01000111",
		6811 => "01110000",
		6812 => "11111001",
		6813 => "11111111",
		6814 => "11111111",
		6815 => "11111111",
		6816 => "11111111",
		6817 => "11111111",
		6818 => "11111111",
		6819 => "11111111",
		6820 => "11111111",
		6821 => "11111111",
		6822 => "11111111",
		6823 => "11001011",
		6824 => "01011110",
		6825 => "01000111",
		6826 => "01010011",
		6827 => "10000111",
		6828 => "11110011",
		6829 => "11010001",
		6830 => "01000111",
		6831 => "01000111",
		6832 => "01000111",
		6833 => "01011001",
		6834 => "11011100",
		6835 => "10000111",
		6836 => "01000111",
		6837 => "01000111",
		6838 => "01101010",
		6839 => "01000111",
		6840 => "10101110",
		6841 => "11111111",
		6842 => "11111111",
		6843 => "11111111",
		6844 => "11111111",
		6845 => "11111111",
		6846 => "11111111",
		6847 => "11111111",
		6848 => "11111111",
		6849 => "11111111",
		6850 => "11111111",
		6851 => "11111111",
		6852 => "11111111",
		6853 => "11111111",
		6854 => "11111111",
		6855 => "11111111",
		6856 => "01101010",
		6857 => "01010011",
		6858 => "11011100",
		6859 => "01110101",
		6860 => "01000111",
		6861 => "11100010",
		6862 => "11100010",
		6863 => "01011001",
		6864 => "01000111",
		6865 => "01000111",
		6866 => "01100100",
		6867 => "11111111",
		6868 => "11111111",
		6869 => "10101001",
		6870 => "01110101",
		6871 => "01010011",
		6872 => "10000001",
		6873 => "11100010",
		6874 => "11111111",
		6875 => "11111111",
		6876 => "11111111",
		6877 => "11111111",
		6878 => "11111111",
		6879 => "11111111",
		6880 => "11111111",
		6881 => "11011100",
		6882 => "11101000",
		6883 => "11111111",
		6884 => "11101000",
		6885 => "01111100",
		6886 => "01000111",
		6887 => "01000111",
		6888 => "11101000",
		6889 => "11111111",
		6890 => "11111111",
		6891 => "11111111",
		6892 => "11111111",
		6893 => "11111111",
		6894 => "11111111",
		6895 => "11110011",
		6896 => "01000111",
		6897 => "11111111",
		6898 => "11111111",
		6899 => "11111111",
		6900 => "11111111",
		6901 => "11111111",
		6902 => "11111111",
		6903 => "11111111",
		6904 => "11111111",
		6905 => "11110011",
		6906 => "10000111",
		6907 => "01000111",
		6908 => "11101000",
		6909 => "11111111",
		6910 => "11111111",
		6911 => "11111111",
		6912 => "11111111",
		6913 => "11111111",
		6914 => "11111111",
		6915 => "11111111",
		6916 => "11100010",
		6917 => "11101110",
		6918 => "11111111",
		6919 => "11111111",
		6920 => "11111111",
		6921 => "11111111",
		6922 => "11111111",
		6923 => "11111111",
		6924 => "11111111",
		6925 => "11111111",
		6926 => "11111111",
		6927 => "11101000",
		6928 => "01101010",
		6929 => "11111111",
		6930 => "11111111",
		6931 => "11111111",
		6932 => "11111111",
		6933 => "11111111",
		6934 => "11111111",
		6935 => "11111111",
		6936 => "10111010",
		6937 => "01000111",
		6938 => "11011100",
		6939 => "11010111",
		6940 => "10010011",
		6941 => "01011110",
		6942 => "01110101",
		6943 => "01001101",
		6944 => "10000001",
		6945 => "11111111",
		6946 => "11111111",
		6947 => "11010001",
		6948 => "01000111",
		6949 => "01010011",
		6950 => "11111111",
		6951 => "11111111",
		6952 => "11111111",
		6953 => "11111111",
		6954 => "11111111",
		6955 => "11101110",
		6956 => "11001011",
		6957 => "11001011",
		6958 => "01000111",
		6959 => "10011110",
		6960 => "01000111",
		6961 => "10011110",
		6962 => "10111010",
		6963 => "01001101",
		6964 => "01000111",
		6965 => "01100100",
		6966 => "01110101",
		6967 => "11010001",
		6968 => "11111111",
		6969 => "11111111",
		6970 => "11111111",
		6971 => "11111111",
		6972 => "11111111",
		6973 => "11111111",
		6974 => "11111111",
		6975 => "11111111",
		6976 => "11111111",
		6977 => "11111111",
		6978 => "11111111",
		6979 => "11111111",
		6980 => "11111111",
		6981 => "11111111",
		6982 => "11111111",
		6983 => "11111111",
		6984 => "11111111",
		6985 => "10011110",
		6986 => "01101010",
		6987 => "01001101",
		6988 => "01000111",
		6989 => "01110000",
		6990 => "10111010",
		6991 => "01101010",
		6992 => "01101010",
		6993 => "01111100",
		6994 => "01100100",
		6995 => "11110011",
		6996 => "11010111",
		6997 => "11011100",
		6998 => "11111111",
		6999 => "11111111",
		7000 => "11111111",
		7001 => "11111111",
		7002 => "11101110",
		7003 => "01001101",
		7004 => "01000111",
		7005 => "10110100",
		7006 => "11111111",
		7007 => "11101110",
		7008 => "01101010",
		7009 => "01011110",
		7010 => "10011110",
		7011 => "01111100",
		7012 => "10101001",
		7013 => "11100010",
		7014 => "11110011",
		7015 => "01000111",
		7016 => "10100011",
		7017 => "11111111",
		7018 => "11111111",
		7019 => "11111111",
		7020 => "11111111",
		7021 => "11111111",
		7022 => "11111111",
		7023 => "11111111",
		7024 => "11101000",
		7025 => "11111111",
		7026 => "11111111",
		7027 => "11111111",
		7028 => "11111111",
		7029 => "11111111",
		7030 => "11111111",
		7031 => "11111111",
		7032 => "11111111",
		7033 => "11111111",
		7034 => "11111111",
		7035 => "11111111",
		7036 => "11111111",
		7037 => "11111111",
		7038 => "11111111",
		7039 => "11111111",
		7040 => "11111111",
		7041 => "11111111",
		7042 => "11111111",
		7043 => "11111111",
		7044 => "10101110",
		7045 => "10111010",
		7046 => "11111111",
		7047 => "11111111",
		7048 => "11111111",
		7049 => "11111111",
		7050 => "11111111",
		7051 => "11111111",
		7052 => "11111111",
		7053 => "11111111",
		7054 => "11111111",
		7055 => "11000101",
		7056 => "10000001",
		7057 => "11111111",
		7058 => "11111111",
		7059 => "11111111",
		7060 => "11111111",
		7061 => "11111111",
		7062 => "11111111",
		7063 => "11111111",
		7064 => "10100011",
		7065 => "01000111",
		7066 => "11111001",
		7067 => "11111111",
		7068 => "11111111",
		7069 => "11111111",
		7070 => "11111111",
		7071 => "11000101",
		7072 => "01000111",
		7073 => "10011110",
		7074 => "10000111",
		7075 => "01001101",
		7076 => "01010011",
		7077 => "01000111",
		7078 => "10110100",
		7079 => "11111111",
		7080 => "11111111",
		7081 => "11111111",
		7082 => "10111010",
		7083 => "01001101",
		7084 => "01000111",
		7085 => "01010011",
		7086 => "01001101",
		7087 => "01100100",
		7088 => "01011001",
		7089 => "11111001",
		7090 => "11011100",
		7091 => "01000111",
		7092 => "01000111",
		7093 => "11001011",
		7094 => "11111111",
		7095 => "11111111",
		7096 => "11111111",
		7097 => "11111111",
		7098 => "11111111",
		7099 => "11111111",
		7100 => "11111111",
		7101 => "11111111",
		7102 => "11111111",
		7103 => "11111111",
		7104 => "11111111",
		7105 => "11111111",
		7106 => "11111111",
		7107 => "11111111",
		7108 => "11111111",
		7109 => "11111111",
		7110 => "11111111",
		7111 => "11111111",
		7112 => "11111111",
		7113 => "11111111",
		7114 => "11111111",
		7115 => "10011000",
		7116 => "01000111",
		7117 => "01111100",
		7118 => "11111111",
		7119 => "11000101",
		7120 => "01000111",
		7121 => "01111100",
		7122 => "01000111",
		7123 => "01011001",
		7124 => "01000111",
		7125 => "01000111",
		7126 => "10001100",
		7127 => "11111111",
		7128 => "11111111",
		7129 => "11111111",
		7130 => "10001100",
		7131 => "01000111",
		7132 => "01011110",
		7133 => "01000111",
		7134 => "01110101",
		7135 => "01000111",
		7136 => "01001101",
		7137 => "11011100",
		7138 => "11111111",
		7139 => "11111111",
		7140 => "11111111",
		7141 => "11111111",
		7142 => "11111111",
		7143 => "01011001",
		7144 => "10001100",
		7145 => "11111111",
		7146 => "11111111",
		7147 => "11111111",
		7148 => "11111111",
		7149 => "11111111",
		7150 => "11111111",
		7151 => "11111111",
		7152 => "11111111",
		7153 => "11111111",
		7154 => "11111111",
		7155 => "11111111",
		7156 => "11111111",
		7157 => "11111111",
		7158 => "11111111",
		7159 => "11111111",
		7160 => "11111111",
		7161 => "11111111",
		7162 => "11111111",
		7163 => "11111111",
		7164 => "11111111",
		7165 => "11111111",
		7166 => "11111111",
		7167 => "11111111",
		7168 => "11111111",
		7169 => "11111111",
		7170 => "11111111",
		7171 => "11111111",
		7172 => "10000111",
		7173 => "01011110",
		7174 => "10011000",
		7175 => "10110100",
		7176 => "11010001",
		7177 => "11111111",
		7178 => "11111111",
		7179 => "11111111",
		7180 => "11111111",
		7181 => "11111111",
		7182 => "11111111",
		7183 => "01111100",
		7184 => "10110100",
		7185 => "11111111",
		7186 => "11111111",
		7187 => "11111111",
		7188 => "11111111",
		7189 => "11111111",
		7190 => "11111111",
		7191 => "11111111",
		7192 => "10001100",
		7193 => "01011110",
		7194 => "11111111",
		7195 => "11111111",
		7196 => "11111111",
		7197 => "11111111",
		7198 => "11111111",
		7199 => "11111111",
		7200 => "11000101",
		7201 => "01010011",
		7202 => "01100100",
		7203 => "10010011",
		7204 => "11110011",
		7205 => "10011110",
		7206 => "01000111",
		7207 => "10010011",
		7208 => "10100011",
		7209 => "10000111",
		7210 => "01000111",
		7211 => "01000111",
		7212 => "01000111",
		7213 => "10001100",
		7214 => "10000111",
		7215 => "01000111",
		7216 => "10100011",
		7217 => "11111111",
		7218 => "11111111",
		7219 => "10000111",
		7220 => "01000111",
		7221 => "10001100",
		7222 => "11111111",
		7223 => "11111111",
		7224 => "11111111",
		7225 => "11111111",
		7226 => "11111111",
		7227 => "11111111",
		7228 => "11111111",
		7229 => "11111111",
		7230 => "11111111",
		7231 => "11111111",
		7232 => "11111111",
		7233 => "11111111",
		7234 => "11111111",
		7235 => "11111111",
		7236 => "11111111",
		7237 => "11111111",
		7238 => "11111111",
		7239 => "11111111",
		7240 => "11111111",
		7241 => "11111111",
		7242 => "11101110",
		7243 => "01000111",
		7244 => "01000111",
		7245 => "10111010",
		7246 => "11111111",
		7247 => "11111111",
		7248 => "01011001",
		7249 => "01011001",
		7250 => "10011110",
		7251 => "01110000",
		7252 => "01000111",
		7253 => "01011110",
		7254 => "01000111",
		7255 => "01100100",
		7256 => "10000111",
		7257 => "01011001",
		7258 => "01000111",
		7259 => "10100011",
		7260 => "11111111",
		7261 => "10110100",
		7262 => "01110101",
		7263 => "10011110",
		7264 => "11100010",
		7265 => "11111111",
		7266 => "11111111",
		7267 => "11111111",
		7268 => "11111111",
		7269 => "11111111",
		7270 => "11111111",
		7271 => "01110000",
		7272 => "01110000",
		7273 => "11111111",
		7274 => "11111111",
		7275 => "11111111",
		7276 => "11111111",
		7277 => "11111111",
		7278 => "11111111",
		7279 => "11111111",
		7280 => "11111111",
		7281 => "10101001",
		7282 => "11111111",
		7283 => "11111111",
		7284 => "11111111",
		7285 => "11111111",
		7286 => "11111111",
		7287 => "11111111",
		7288 => "11111111",
		7289 => "11111111",
		7290 => "11111111",
		7291 => "11111111",
		7292 => "11111111",
		7293 => "11111111",
		7294 => "11111111",
		7295 => "11111111",
		7296 => "11111111",
		7297 => "11111111",
		7298 => "11111111",
		7299 => "11111111",
		7300 => "01101010",
		7301 => "01000111",
		7302 => "01000111",
		7303 => "01000111",
		7304 => "01000111",
		7305 => "01000111",
		7306 => "01101010",
		7307 => "10000111",
		7308 => "10100011",
		7309 => "11000000",
		7310 => "01111100",
		7311 => "01001101",
		7312 => "11101110",
		7313 => "11111111",
		7314 => "11111111",
		7315 => "11111111",
		7316 => "11111111",
		7317 => "11111111",
		7318 => "11111111",
		7319 => "11111111",
		7320 => "01110101",
		7321 => "01111100",
		7322 => "11111111",
		7323 => "11111111",
		7324 => "11111111",
		7325 => "11111111",
		7326 => "11111111",
		7327 => "11111111",
		7328 => "11111111",
		7329 => "11111111",
		7330 => "11111111",
		7331 => "11111111",
		7332 => "11111111",
		7333 => "11111111",
		7334 => "10101001",
		7335 => "01101010",
		7336 => "01000111",
		7337 => "01000111",
		7338 => "10011000",
		7339 => "10010011",
		7340 => "01000111",
		7341 => "01000111",
		7342 => "01000111",
		7343 => "01000111",
		7344 => "10010011",
		7345 => "11110011",
		7346 => "10100011",
		7347 => "10100011",
		7348 => "01001101",
		7349 => "10100011",
		7350 => "11111111",
		7351 => "10101001",
		7352 => "10100011",
		7353 => "10100011",
		7354 => "10100011",
		7355 => "11000101",
		7356 => "11111111",
		7357 => "11111111",
		7358 => "11111111",
		7359 => "11111111",
		7360 => "11111111",
		7361 => "11111111",
		7362 => "11111111",
		7363 => "11111111",
		7364 => "11111111",
		7365 => "11111001",
		7366 => "10110100",
		7367 => "10000111",
		7368 => "01110101",
		7369 => "10100011",
		7370 => "11111111",
		7371 => "01011110",
		7372 => "01110000",
		7373 => "10100011",
		7374 => "11000000",
		7375 => "11111001",
		7376 => "01000111",
		7377 => "01000111",
		7378 => "01000111",
		7379 => "01000111",
		7380 => "01000111",
		7381 => "11011100",
		7382 => "11001011",
		7383 => "01111100",
		7384 => "01011110",
		7385 => "10000111",
		7386 => "11000000",
		7387 => "11111111",
		7388 => "11111111",
		7389 => "11111111",
		7390 => "11111111",
		7391 => "11111111",
		7392 => "11111111",
		7393 => "11111111",
		7394 => "11111111",
		7395 => "11111111",
		7396 => "11111111",
		7397 => "11111111",
		7398 => "11111111",
		7399 => "10001100",
		7400 => "01011001",
		7401 => "11111111",
		7402 => "11111111",
		7403 => "11111111",
		7404 => "11111111",
		7405 => "11111111",
		7406 => "11111111",
		7407 => "11111111",
		7408 => "11111111",
		7409 => "01110101",
		7410 => "10111010",
		7411 => "11111111",
		7412 => "11111111",
		7413 => "11111111",
		7414 => "11111111",
		7415 => "11111111",
		7416 => "11111111",
		7417 => "11111111",
		7418 => "11111111",
		7419 => "11111111",
		7420 => "11111111",
		7421 => "11111111",
		7422 => "11111111",
		7423 => "11111111",
		7424 => "11111111",
		7425 => "11111111",
		7426 => "11111111",
		7427 => "11111001",
		7428 => "01011110",
		7429 => "11110011",
		7430 => "11010001",
		7431 => "10101110",
		7432 => "10010011",
		7433 => "01110101",
		7434 => "01000111",
		7435 => "01000111",
		7436 => "01000111",
		7437 => "01000111",
		7438 => "01000111",
		7439 => "11000000",
		7440 => "11111111",
		7441 => "11111111",
		7442 => "11111111",
		7443 => "11111111",
		7444 => "11111111",
		7445 => "11111111",
		7446 => "11111111",
		7447 => "11111111",
		7448 => "01011110",
		7449 => "10010011",
		7450 => "11111111",
		7451 => "11111111",
		7452 => "11111111",
		7453 => "11111111",
		7454 => "11111111",
		7455 => "11111111",
		7456 => "11111111",
		7457 => "11111111",
		7458 => "11111111",
		7459 => "11111111",
		7460 => "11111111",
		7461 => "11111111",
		7462 => "11111111",
		7463 => "11111111",
		7464 => "11111111",
		7465 => "11000000",
		7466 => "11000000",
		7467 => "11111111",
		7468 => "11001011",
		7469 => "01000111",
		7470 => "01101010",
		7471 => "01011110",
		7472 => "01111100",
		7473 => "10100011",
		7474 => "01000111",
		7475 => "01000111",
		7476 => "01000111",
		7477 => "10010011",
		7478 => "11111111",
		7479 => "11111111",
		7480 => "11111111",
		7481 => "11111111",
		7482 => "11111001",
		7483 => "11000000",
		7484 => "11000101",
		7485 => "11111111",
		7486 => "11111111",
		7487 => "11111111",
		7488 => "11111111",
		7489 => "11111111",
		7490 => "11111111",
		7491 => "11111111",
		7492 => "11111111",
		7493 => "10011110",
		7494 => "11010111",
		7495 => "11111111",
		7496 => "11111111",
		7497 => "11111001",
		7498 => "11111111",
		7499 => "10010011",
		7500 => "01000111",
		7501 => "01000111",
		7502 => "01000111",
		7503 => "11010001",
		7504 => "01000111",
		7505 => "01110000",
		7506 => "01000111",
		7507 => "01110101",
		7508 => "11100010",
		7509 => "11111111",
		7510 => "10110100",
		7511 => "10011110",
		7512 => "11111111",
		7513 => "11111111",
		7514 => "11111111",
		7515 => "11111111",
		7516 => "11110011",
		7517 => "11111111",
		7518 => "11111111",
		7519 => "11111111",
		7520 => "11111111",
		7521 => "11111111",
		7522 => "11111111",
		7523 => "11111111",
		7524 => "11111111",
		7525 => "11111111",
		7526 => "11111111",
		7527 => "10100011",
		7528 => "01000111",
		7529 => "11111001",
		7530 => "11111111",
		7531 => "11111111",
		7532 => "11111111",
		7533 => "11111111",
		7534 => "11111111",
		7535 => "11111111",
		7536 => "11111111",
		7537 => "01110101",
		7538 => "01000111",
		7539 => "10011000",
		7540 => "11100010",
		7541 => "11111111",
		7542 => "11111111",
		7543 => "11111111",
		7544 => "11111111",
		7545 => "11111111",
		7546 => "11111111",
		7547 => "11111111",
		7548 => "11111111",
		7549 => "11111111",
		7550 => "11111111",
		7551 => "11111111",
		7552 => "11111111",
		7553 => "11111111",
		7554 => "11111111",
		7555 => "11111001",
		7556 => "11011100",
		7557 => "11111111",
		7558 => "11111111",
		7559 => "11111111",
		7560 => "11111111",
		7561 => "11111111",
		7562 => "11111111",
		7563 => "11100010",
		7564 => "11000101",
		7565 => "10101110",
		7566 => "11101110",
		7567 => "11111111",
		7568 => "11111111",
		7569 => "11111111",
		7570 => "11111111",
		7571 => "11111111",
		7572 => "11111111",
		7573 => "11111111",
		7574 => "11111111",
		7575 => "11111111",
		7576 => "01000111",
		7577 => "01100100",
		7578 => "11111111",
		7579 => "11111111",
		7580 => "11111111",
		7581 => "11111111",
		7582 => "11101000",
		7583 => "10011110",
		7584 => "11111001",
		7585 => "11111111",
		7586 => "11111111",
		7587 => "11101000",
		7588 => "01011110",
		7589 => "11000000",
		7590 => "11111111",
		7591 => "11111111",
		7592 => "11101000",
		7593 => "01001101",
		7594 => "10000001",
		7595 => "11111111",
		7596 => "11111111",
		7597 => "01011110",
		7598 => "01000111",
		7599 => "01000111",
		7600 => "10101001",
		7601 => "01011110",
		7602 => "01110000",
		7603 => "11111111",
		7604 => "01011110",
		7605 => "10001100",
		7606 => "11111111",
		7607 => "11111111",
		7608 => "11111111",
		7609 => "11111111",
		7610 => "11111111",
		7611 => "11111111",
		7612 => "11111111",
		7613 => "11111111",
		7614 => "11111111",
		7615 => "11111111",
		7616 => "11111111",
		7617 => "11111111",
		7618 => "11111111",
		7619 => "11111111",
		7620 => "11111111",
		7621 => "11111111",
		7622 => "11111111",
		7623 => "11111111",
		7624 => "11111111",
		7625 => "11111111",
		7626 => "11111111",
		7627 => "10001100",
		7628 => "01011110",
		7629 => "11010111",
		7630 => "01000111",
		7631 => "10011110",
		7632 => "01111100",
		7633 => "01000111",
		7634 => "01000111",
		7635 => "10101001",
		7636 => "11111111",
		7637 => "11111111",
		7638 => "10011000",
		7639 => "01001101",
		7640 => "11010001",
		7641 => "11111111",
		7642 => "11111111",
		7643 => "10111010",
		7644 => "01000111",
		7645 => "11010111",
		7646 => "11111111",
		7647 => "11111111",
		7648 => "11101110",
		7649 => "01111100",
		7650 => "11010111",
		7651 => "11111111",
		7652 => "11111111",
		7653 => "11111111",
		7654 => "11111111",
		7655 => "10011000",
		7656 => "01000111",
		7657 => "11101000",
		7658 => "11111111",
		7659 => "11111111",
		7660 => "11111111",
		7661 => "11111111",
		7662 => "11111111",
		7663 => "11111111",
		7664 => "11111111",
		7665 => "10001100",
		7666 => "11000000",
		7667 => "10010011",
		7668 => "01011110",
		7669 => "01100100",
		7670 => "10101001",
		7671 => "11101000",
		7672 => "11111111",
		7673 => "11111111",
		7674 => "11111111",
		7675 => "11111111",
		7676 => "11111111",
		7677 => "11111111",
		7678 => "11111111",
		7679 => "11111111",
		7680 => "11111111",
		7681 => "11111111",
		7682 => "11111111",
		7683 => "11111111",
		7684 => "11111111",
		7685 => "11111111",
		7686 => "11111111",
		7687 => "11111111",
		7688 => "11111111",
		7689 => "11111111",
		7690 => "11111111",
		7691 => "11111111",
		7692 => "11111111",
		7693 => "11111111",
		7694 => "11111111",
		7695 => "11111111",
		7696 => "11111111",
		7697 => "11111111",
		7698 => "11111111",
		7699 => "11111111",
		7700 => "11111111",
		7701 => "11111111",
		7702 => "11111111",
		7703 => "11111111",
		7704 => "01000111",
		7705 => "01000111",
		7706 => "11011100",
		7707 => "11111111",
		7708 => "11111111",
		7709 => "11111111",
		7710 => "01110101",
		7711 => "01000111",
		7712 => "10100011",
		7713 => "11111111",
		7714 => "11111111",
		7715 => "10101001",
		7716 => "01000111",
		7717 => "01001101",
		7718 => "10011000",
		7719 => "10011110",
		7720 => "01011110",
		7721 => "01000111",
		7722 => "10001100",
		7723 => "11111111",
		7724 => "11111111",
		7725 => "10001100",
		7726 => "01000111",
		7727 => "01000111",
		7728 => "01000111",
		7729 => "01001101",
		7730 => "11010111",
		7731 => "11111001",
		7732 => "01001101",
		7733 => "10010011",
		7734 => "11111111",
		7735 => "11001011",
		7736 => "01101010",
		7737 => "01000111",
		7738 => "01000111",
		7739 => "10000111",
		7740 => "10010011",
		7741 => "10111010",
		7742 => "11111111",
		7743 => "11111111",
		7744 => "11111111",
		7745 => "11111111",
		7746 => "11111111",
		7747 => "11111111",
		7748 => "11111111",
		7749 => "11011100",
		7750 => "10010011",
		7751 => "01110101",
		7752 => "01110101",
		7753 => "10100011",
		7754 => "11111111",
		7755 => "10011000",
		7756 => "01011001",
		7757 => "11111111",
		7758 => "10001100",
		7759 => "01000111",
		7760 => "01000111",
		7761 => "01000111",
		7762 => "01000111",
		7763 => "11010001",
		7764 => "11111111",
		7765 => "11111111",
		7766 => "10100011",
		7767 => "01000111",
		7768 => "01010011",
		7769 => "10001100",
		7770 => "10000111",
		7771 => "01001101",
		7772 => "01000111",
		7773 => "10011000",
		7774 => "11111111",
		7775 => "11111111",
		7776 => "10011000",
		7777 => "01000111",
		7778 => "01011001",
		7779 => "11111001",
		7780 => "11111111",
		7781 => "11111111",
		7782 => "11101000",
		7783 => "01001101",
		7784 => "01000111",
		7785 => "11101000",
		7786 => "11111111",
		7787 => "11111111",
		7788 => "11111111",
		7789 => "11111111",
		7790 => "11111111",
		7791 => "11111111",
		7792 => "11111111",
		7793 => "11001011",
		7794 => "11111111",
		7795 => "11111111",
		7796 => "11111111",
		7797 => "10011000",
		7798 => "01111100",
		7799 => "01011110",
		7800 => "01101010",
		7801 => "10110100",
		7802 => "11101110",
		7803 => "11111111",
		7804 => "11111111",
		7805 => "11111111",
		7806 => "11111111",
		7807 => "11111111",
		7808 => "11111111",
		7809 => "11111111",
		7810 => "11111111",
		7811 => "11111111",
		7812 => "11111111",
		7813 => "11111111",
		7814 => "11111111",
		7815 => "11111111",
		7816 => "11111111",
		7817 => "11111111",
		7818 => "11111111",
		7819 => "11111111",
		7820 => "11111111",
		7821 => "11111111",
		7822 => "11111111",
		7823 => "11111111",
		7824 => "11111111",
		7825 => "11111111",
		7826 => "11111111",
		7827 => "11111111",
		7828 => "11111111",
		7829 => "11111111",
		7830 => "11111111",
		7831 => "11111111",
		7832 => "01000111",
		7833 => "01000111",
		7834 => "01011110",
		7835 => "11001011",
		7836 => "11100010",
		7837 => "10011000",
		7838 => "01000111",
		7839 => "01000111",
		7840 => "01001101",
		7841 => "11101110",
		7842 => "10101001",
		7843 => "01010011",
		7844 => "01000111",
		7845 => "01011110",
		7846 => "01010011",
		7847 => "01000111",
		7848 => "01111100",
		7849 => "01010011",
		7850 => "10001100",
		7851 => "11111111",
		7852 => "11111111",
		7853 => "11010111",
		7854 => "01000111",
		7855 => "01101010",
		7856 => "01010011",
		7857 => "01110000",
		7858 => "11111111",
		7859 => "10011000",
		7860 => "01000111",
		7861 => "11010111",
		7862 => "11010111",
		7863 => "01101010",
		7864 => "01011110",
		7865 => "01000111",
		7866 => "01011110",
		7867 => "01100100",
		7868 => "01011110",
		7869 => "01010011",
		7870 => "11111111",
		7871 => "11111111",
		7872 => "11111111",
		7873 => "11111111",
		7874 => "11111111",
		7875 => "11111111",
		7876 => "10111010",
		7877 => "01011001",
		7878 => "01011110",
		7879 => "01000111",
		7880 => "01000111",
		7881 => "01010011",
		7882 => "11101110",
		7883 => "10111010",
		7884 => "01000111",
		7885 => "11010001",
		7886 => "11111111",
		7887 => "01100100",
		7888 => "01010011",
		7889 => "01000111",
		7890 => "01011110",
		7891 => "11111001",
		7892 => "11111111",
		7893 => "11111111",
		7894 => "10010011",
		7895 => "01000111",
		7896 => "10010011",
		7897 => "01011110",
		7898 => "01100100",
		7899 => "01110101",
		7900 => "01000111",
		7901 => "01000111",
		7902 => "11000101",
		7903 => "10101110",
		7904 => "01001101",
		7905 => "01000111",
		7906 => "01000111",
		7907 => "01110101",
		7908 => "10111010",
		7909 => "10110100",
		7910 => "01011001",
		7911 => "01000111",
		7912 => "01000111",
		7913 => "11101000",
		7914 => "11111111",
		7915 => "11111111",
		7916 => "11111111",
		7917 => "11111111",
		7918 => "11111111",
		7919 => "11111111",
		7920 => "11111111",
		7921 => "11111111",
		7922 => "11111111",
		7923 => "11111111",
		7924 => "11111111",
		7925 => "10101110",
		7926 => "11000101",
		7927 => "11111111",
		7928 => "11011100",
		7929 => "10100011",
		7930 => "01101010",
		7931 => "01110101",
		7932 => "10111010",
		7933 => "11111111",
		7934 => "11111111",
		7935 => "11111111",
		7936 => "11111111",
		7937 => "11111111",
		7938 => "11111111",
		7939 => "11111111",
		7940 => "11111111",
		7941 => "11111111",
		7942 => "11111111",
		7943 => "11111111",
		7944 => "11111111",
		7945 => "11111111",
		7946 => "11111111",
		7947 => "11111111",
		7948 => "11111111",
		7949 => "11111111",
		7950 => "11111111",
		7951 => "11111111",
		7952 => "11111111",
		7953 => "11111111",
		7954 => "11111111",
		7955 => "11111111",
		7956 => "11111111",
		7957 => "11111111",
		7958 => "11111111",
		7959 => "11111111",
		7960 => "01000111",
		7961 => "10011000",
		7962 => "01011110",
		7963 => "01000111",
		7964 => "01000111",
		7965 => "01000111",
		7966 => "01110000",
		7967 => "01000111",
		7968 => "01010011",
		7969 => "01000111",
		7970 => "01000111",
		7971 => "01101010",
		7972 => "01000111",
		7973 => "10011110",
		7974 => "11111111",
		7975 => "11111111",
		7976 => "11111111",
		7977 => "01101010",
		7978 => "10000111",
		7979 => "11111111",
		7980 => "11010001",
		7981 => "10001100",
		7982 => "01111100",
		7983 => "01011001",
		7984 => "01000111",
		7985 => "10010011",
		7986 => "11001011",
		7987 => "01000111",
		7988 => "10010011",
		7989 => "11111111",
		7990 => "10011110",
		7991 => "10111010",
		7992 => "01101010",
		7993 => "01000111",
		7994 => "01000111",
		7995 => "10000111",
		7996 => "11000101",
		7997 => "01000111",
		7998 => "11010111",
		7999 => "11111111",
		8000 => "11111111",
		8001 => "11111111",
		8002 => "11111111",
		8003 => "11110011",
		8004 => "01001101",
		8005 => "10110100",
		8006 => "01101010",
		8007 => "01000111",
		8008 => "01011001",
		8009 => "01110000",
		8010 => "10101001",
		8011 => "11111111",
		8012 => "01110000",
		8013 => "01010011",
		8014 => "11101110",
		8015 => "10011000",
		8016 => "01000111",
		8017 => "01000111",
		8018 => "10100011",
		8019 => "10000111",
		8020 => "11111001",
		8021 => "11111111",
		8022 => "10001100",
		8023 => "01001101",
		8024 => "11111111",
		8025 => "11111111",
		8026 => "11111111",
		8027 => "10101110",
		8028 => "01000111",
		8029 => "10000001",
		8030 => "01000111",
		8031 => "01000111",
		8032 => "01111100",
		8033 => "01000111",
		8034 => "01110000",
		8035 => "01010011",
		8036 => "01000111",
		8037 => "01000111",
		8038 => "01110101",
		8039 => "10011000",
		8040 => "01000111",
		8041 => "11101000",
		8042 => "11111111",
		8043 => "11111111",
		8044 => "11111111",
		8045 => "11111111",
		8046 => "11111111",
		8047 => "11111111",
		8048 => "11111111",
		8049 => "11111111",
		8050 => "11111111",
		8051 => "11111111",
		8052 => "11111111",
		8053 => "10111010",
		8054 => "10111010",
		8055 => "11111111",
		8056 => "11110011",
		8057 => "10110100",
		8058 => "01110101",
		8059 => "01000111",
		8060 => "01000111",
		8061 => "11111111",
		8062 => "11111111",
		8063 => "11111111",
		8064 => "11111111",
		8065 => "11111111",
		8066 => "11111111",
		8067 => "11111111",
		8068 => "11111111",
		8069 => "11111111",
		8070 => "11111111",
		8071 => "11111111",
		8072 => "11111111",
		8073 => "11111111",
		8074 => "11111111",
		8075 => "11101000",
		8076 => "10110100",
		8077 => "11010111",
		8078 => "11111111",
		8079 => "11111111",
		8080 => "11111111",
		8081 => "11111111",
		8082 => "11111111",
		8083 => "11111111",
		8084 => "11111111",
		8085 => "11111111",
		8086 => "11111111",
		8087 => "11111111",
		8088 => "01000111",
		8089 => "10111010",
		8090 => "11111111",
		8091 => "11011100",
		8092 => "10110100",
		8093 => "11100010",
		8094 => "11010001",
		8095 => "01000111",
		8096 => "11000000",
		8097 => "10100011",
		8098 => "11010001",
		8099 => "11111111",
		8100 => "01010011",
		8101 => "10000111",
		8102 => "11111111",
		8103 => "11111111",
		8104 => "11111111",
		8105 => "01110101",
		8106 => "01110101",
		8107 => "11111111",
		8108 => "01110101",
		8109 => "01000111",
		8110 => "01000111",
		8111 => "01011001",
		8112 => "01000111",
		8113 => "10100011",
		8114 => "10010011",
		8115 => "01001101",
		8116 => "11111001",
		8117 => "11111111",
		8118 => "11111001",
		8119 => "10100011",
		8120 => "01110000",
		8121 => "01000111",
		8122 => "01000111",
		8123 => "10000111",
		8124 => "10010011",
		8125 => "01001101",
		8126 => "11101000",
		8127 => "11111111",
		8128 => "11111111",
		8129 => "11111111",
		8130 => "11111111",
		8131 => "11110011",
		8132 => "01110101",
		8133 => "10011000",
		8134 => "01100100",
		8135 => "01000111",
		8136 => "01000111",
		8137 => "10011000",
		8138 => "11011100",
		8139 => "11111111",
		8140 => "11100010",
		8141 => "01000111",
		8142 => "10011110",
		8143 => "10110100",
		8144 => "01000111",
		8145 => "01000111",
		8146 => "01000111",
		8147 => "01000111",
		8148 => "11000101",
		8149 => "11111111",
		8150 => "10001100",
		8151 => "01011110",
		8152 => "11111111",
		8153 => "11111111",
		8154 => "11111111",
		8155 => "10011110",
		8156 => "01001101",
		8157 => "11111111",
		8158 => "11010001",
		8159 => "11100010",
		8160 => "11101000",
		8161 => "01000111",
		8162 => "10110100",
		8163 => "11111111",
		8164 => "11010001",
		8165 => "11110011",
		8166 => "11111111",
		8167 => "10111010",
		8168 => "01000111",
		8169 => "11101000",
		8170 => "11111111",
		8171 => "11111111",
		8172 => "11111111",
		8173 => "11111111",
		8174 => "11111111",
		8175 => "11111111",
		8176 => "11111111",
		8177 => "11111111",
		8178 => "11111111",
		8179 => "11111111",
		8180 => "11111111",
		8181 => "10111010",
		8182 => "10011000",
		8183 => "10001100",
		8184 => "01001101",
		8185 => "01000111",
		8186 => "01000111",
		8187 => "10000111",
		8188 => "11001011",
		8189 => "11111111",
		8190 => "11111111",
		8191 => "11111111",
		8192 => "11111111",
		8193 => "11111111",
		8194 => "11111111",
		8195 => "11111111",
		8196 => "01011001",
		8197 => "01000111",
		8198 => "01110101",
		8199 => "11111111",
		8200 => "11111111",
		8201 => "11111111",
		8202 => "11000000",
		8203 => "01000111",
		8204 => "01000111",
		8205 => "01000111",
		8206 => "10011000",
		8207 => "11111111",
		8208 => "11111111",
		8209 => "11111111",
		8210 => "11111111",
		8211 => "11111111",
		8212 => "11111111",
		8213 => "11111111",
		8214 => "11111111",
		8215 => "11111111",
		8216 => "01000111",
		8217 => "10111010",
		8218 => "11111111",
		8219 => "11111111",
		8220 => "11111111",
		8221 => "11111111",
		8222 => "11100010",
		8223 => "01000111",
		8224 => "10111010",
		8225 => "11111111",
		8226 => "11111111",
		8227 => "11111111",
		8228 => "01110000",
		8229 => "01110000",
		8230 => "11111111",
		8231 => "11111111",
		8232 => "11111111",
		8233 => "10000001",
		8234 => "01100100",
		8235 => "11111111",
		8236 => "01100100",
		8237 => "01001101",
		8238 => "10000001",
		8239 => "11101000",
		8240 => "01001101",
		8241 => "10010011",
		8242 => "10001100",
		8243 => "01010011",
		8244 => "10101110",
		8245 => "11111111",
		8246 => "11111111",
		8247 => "11111111",
		8248 => "11111111",
		8249 => "11111111",
		8250 => "10011110",
		8251 => "10011110",
		8252 => "01101010",
		8253 => "11001011",
		8254 => "11111111",
		8255 => "11111111",
		8256 => "11111111",
		8257 => "11111111",
		8258 => "11111111",
		8259 => "11111111",
		8260 => "11011100",
		8261 => "10100011",
		8262 => "10001010",
		8263 => "10100001",
		8264 => "11010001",
		8265 => "11010001",
		8266 => "11111111",
		8267 => "11111111",
		8268 => "11111111",
		8269 => "01101010",
		8270 => "01111100",
		8271 => "10101110",
		8272 => "01000111",
		8273 => "10010011",
		8274 => "01100100",
		8275 => "01000111",
		8276 => "10101001",
		8277 => "11111111",
		8278 => "01111100",
		8279 => "01011110",
		8280 => "11111111",
		8281 => "11111111",
		8282 => "11111111",
		8283 => "10000111",
		8284 => "01100100",
		8285 => "11111111",
		8286 => "11111111",
		8287 => "11111111",
		8288 => "11011100",
		8289 => "01000111",
		8290 => "11000000",
		8291 => "11111111",
		8292 => "11111111",
		8293 => "11111111",
		8294 => "11111111",
		8295 => "10111010",
		8296 => "01000111",
		8297 => "11101000",
		8298 => "11111111",
		8299 => "11111111",
		8300 => "11111111",
		8301 => "11111111",
		8302 => "11111111",
		8303 => "11111111",
		8304 => "11111111",
		8305 => "11001011",
		8306 => "11011100",
		8307 => "11110011",
		8308 => "10110100",
		8309 => "01100100",
		8310 => "01000111",
		8311 => "01000111",
		8312 => "01011110",
		8313 => "10101001",
		8314 => "11101110",
		8315 => "11111111",
		8316 => "11111111",
		8317 => "11111111",
		8318 => "11111111",
		8319 => "11111111",
		8320 => "11111111",
		8321 => "11111111",
		8322 => "11111111",
		8323 => "11110011",
		8324 => "01101010",
		8325 => "11001011",
		8326 => "11111111",
		8327 => "11111111",
		8328 => "11111111",
		8329 => "11101000",
		8330 => "01001101",
		8331 => "01000111",
		8332 => "10000111",
		8333 => "10001100",
		8334 => "01001101",
		8335 => "11011100",
		8336 => "11111111",
		8337 => "11111111",
		8338 => "11111111",
		8339 => "11111111",
		8340 => "11111111",
		8341 => "11111111",
		8342 => "11111111",
		8343 => "11111111",
		8344 => "01000111",
		8345 => "10110100",
		8346 => "11111111",
		8347 => "11111111",
		8348 => "11111111",
		8349 => "11111111",
		8350 => "11101000",
		8351 => "01000111",
		8352 => "10101001",
		8353 => "11111111",
		8354 => "11111111",
		8355 => "11111111",
		8356 => "10010011",
		8357 => "01011001",
		8358 => "11111111",
		8359 => "11111111",
		8360 => "11111111",
		8361 => "10010011",
		8362 => "01010011",
		8363 => "11111111",
		8364 => "10011000",
		8365 => "01000111",
		8366 => "01111100",
		8367 => "11101000",
		8368 => "10000001",
		8369 => "01001101",
		8370 => "11000000",
		8371 => "01001101",
		8372 => "01000111",
		8373 => "11101000",
		8374 => "11111111",
		8375 => "11111111",
		8376 => "11111111",
		8377 => "11111111",
		8378 => "11111111",
		8379 => "11111111",
		8380 => "11111111",
		8381 => "11111111",
		8382 => "11111111",
		8383 => "11111111",
		8384 => "11111111",
		8385 => "11111111",
		8386 => "11111111",
		8387 => "11111111",
		8388 => "11111111",
		8389 => "11111111",
		8390 => "11111111",
		8391 => "11111111",
		8392 => "11111111",
		8393 => "11111111",
		8394 => "11111111",
		8395 => "11101110",
		8396 => "01001101",
		8397 => "01000111",
		8398 => "10100011",
		8399 => "01101010",
		8400 => "01101010",
		8401 => "10111010",
		8402 => "01011001",
		8403 => "01001101",
		8404 => "11011100",
		8405 => "11111111",
		8406 => "01100100",
		8407 => "01110000",
		8408 => "11111111",
		8409 => "11111111",
		8410 => "11111111",
		8411 => "01110000",
		8412 => "10000001",
		8413 => "11111111",
		8414 => "11111111",
		8415 => "11111111",
		8416 => "11010001",
		8417 => "01000111",
		8418 => "11010001",
		8419 => "11111111",
		8420 => "11111111",
		8421 => "11111111",
		8422 => "11111111",
		8423 => "10111010",
		8424 => "01000111",
		8425 => "11101000",
		8426 => "11111111",
		8427 => "11111111",
		8428 => "11111111",
		8429 => "11111111",
		8430 => "11111111",
		8431 => "11111111",
		8432 => "11111111",
		8433 => "10111010",
		8434 => "01110000",
		8435 => "01001101",
		8436 => "01000111",
		8437 => "01000111",
		8438 => "01111100",
		8439 => "11000101",
		8440 => "11111111",
		8441 => "11111111",
		8442 => "11111111",
		8443 => "11111111",
		8444 => "11111111",
		8445 => "11111111",
		8446 => "11111111",
		8447 => "11111111",
		8448 => "11111111",
		8449 => "11111111",
		8450 => "11111111",
		8451 => "11100100",
		8452 => "10001100",
		8453 => "11111111",
		8454 => "11111111",
		8455 => "11111111",
		8456 => "11111111",
		8457 => "10000001",
		8458 => "01000111",
		8459 => "01110101",
		8460 => "11111111",
		8461 => "11111111",
		8462 => "10000001",
		8463 => "10101001",
		8464 => "11111111",
		8465 => "11111111",
		8466 => "11111111",
		8467 => "11111111",
		8468 => "11111111",
		8469 => "11111111",
		8470 => "11111111",
		8471 => "11111111",
		8472 => "01000111",
		8473 => "10100011",
		8474 => "11111111",
		8475 => "11111111",
		8476 => "11111111",
		8477 => "11111111",
		8478 => "11111001",
		8479 => "01000111",
		8480 => "10100011",
		8481 => "11111111",
		8482 => "11111111",
		8483 => "11111111",
		8484 => "10101001",
		8485 => "01000111",
		8486 => "11101000",
		8487 => "11111111",
		8488 => "11111111",
		8489 => "10101001",
		8490 => "01000111",
		8491 => "11111001",
		8492 => "11111001",
		8493 => "10101110",
		8494 => "01010011",
		8495 => "01110101",
		8496 => "11001011",
		8497 => "01000111",
		8498 => "01100100",
		8499 => "01011110",
		8500 => "01101010",
		8501 => "11111111",
		8502 => "11111111",
		8503 => "11111111",
		8504 => "11111111",
		8505 => "11111111",
		8506 => "11111111",
		8507 => "11111111",
		8508 => "11111111",
		8509 => "11111111",
		8510 => "11111111",
		8511 => "11111111",
		8512 => "11111111",
		8513 => "11111111",
		8514 => "11111111",
		8515 => "11111111",
		8516 => "11111111",
		8517 => "11111111",
		8518 => "11111111",
		8519 => "11111111",
		8520 => "11111111",
		8521 => "11111111",
		8522 => "11111111",
		8523 => "11111001",
		8524 => "01011001",
		8525 => "01011110",
		8526 => "10100011",
		8527 => "01000111",
		8528 => "10011110",
		8529 => "01000111",
		8530 => "01101010",
		8531 => "11001011",
		8532 => "11111111",
		8533 => "11111111",
		8534 => "01001101",
		8535 => "10001100",
		8536 => "11111111",
		8537 => "11111111",
		8538 => "11111111",
		8539 => "01001101",
		8540 => "10011000",
		8541 => "11111111",
		8542 => "11111111",
		8543 => "11111111",
		8544 => "10111010",
		8545 => "01000111",
		8546 => "11100010",
		8547 => "11111111",
		8548 => "11111111",
		8549 => "11111111",
		8550 => "11111111",
		8551 => "10101001",
		8552 => "01000111",
		8553 => "11111001",
		8554 => "11111111",
		8555 => "11111111",
		8556 => "11111111",
		8557 => "11111111",
		8558 => "11111111",
		8559 => "11111111",
		8560 => "11111111",
		8561 => "11000000",
		8562 => "01000111",
		8563 => "01011001",
		8564 => "10011110",
		8565 => "11101000",
		8566 => "11111111",
		8567 => "11111111",
		8568 => "11111111",
		8569 => "11111111",
		8570 => "11111111",
		8571 => "11111111",
		8572 => "11111111",
		8573 => "11111111",
		8574 => "11111111",
		8575 => "11111111",
		8576 => "11111111",
		8577 => "11111111",
		8578 => "11111111",
		8579 => "11011010",
		8580 => "01111100",
		8581 => "11111111",
		8582 => "11111111",
		8583 => "11111111",
		8584 => "11000101",
		8585 => "01000111",
		8586 => "01001101",
		8587 => "11101000",
		8588 => "11111111",
		8589 => "11111111",
		8590 => "10101110",
		8591 => "10010011",
		8592 => "11111111",
		8593 => "11111111",
		8594 => "11111111",
		8595 => "11111111",
		8596 => "11111111",
		8597 => "11111111",
		8598 => "11111111",
		8599 => "11111111",
		8600 => "01011110",
		8601 => "10001100",
		8602 => "11111111",
		8603 => "11111111",
		8604 => "11111111",
		8605 => "11111111",
		8606 => "11111111",
		8607 => "01000111",
		8608 => "10001100",
		8609 => "11111111",
		8610 => "11111111",
		8611 => "11111111",
		8612 => "11010001",
		8613 => "01000111",
		8614 => "11000101",
		8615 => "11111111",
		8616 => "11111111",
		8617 => "11000000",
		8618 => "01000111",
		8619 => "11011100",
		8620 => "11111111",
		8621 => "11111111",
		8622 => "10101110",
		8623 => "01000111",
		8624 => "01000111",
		8625 => "01010011",
		8626 => "01110000",
		8627 => "01000111",
		8628 => "10110100",
		8629 => "11111111",
		8630 => "11111111",
		8631 => "11111111",
		8632 => "11111111",
		8633 => "11111111",
		8634 => "11111111",
		8635 => "11111111",
		8636 => "11111111",
		8637 => "11111001",
		8638 => "10110100",
		8639 => "11111111",
		8640 => "11111111",
		8641 => "11111111",
		8642 => "11111111",
		8643 => "11111111",
		8644 => "11111111",
		8645 => "11111111",
		8646 => "11111111",
		8647 => "11111111",
		8648 => "11111111",
		8649 => "11111111",
		8650 => "11111111",
		8651 => "11111111",
		8652 => "10101110",
		8653 => "01000111",
		8654 => "01000111",
		8655 => "01000111",
		8656 => "01011001",
		8657 => "01001101",
		8658 => "11101110",
		8659 => "11111111",
		8660 => "11111111",
		8661 => "11101000",
		8662 => "01000111",
		8663 => "10101001",
		8664 => "11111111",
		8665 => "11111111",
		8666 => "11011100",
		8667 => "01000111",
		8668 => "10111010",
		8669 => "11111111",
		8670 => "11111111",
		8671 => "11111111",
		8672 => "10101001",
		8673 => "01000111",
		8674 => "11101110",
		8675 => "11111111",
		8676 => "11111111",
		8677 => "11111111",
		8678 => "11111111",
		8679 => "10011000",
		8680 => "01001101",
		8681 => "11111111",
		8682 => "11111111",
		8683 => "11111111",
		8684 => "11111111",
		8685 => "11111111",
		8686 => "11111111",
		8687 => "11111111",
		8688 => "11111111",
		8689 => "11010001",
		8690 => "01011001",
		8691 => "11111111",
		8692 => "11111111",
		8693 => "11111111",
		8694 => "11111111",
		8695 => "11111111",
		8696 => "11111111",
		8697 => "11111111",
		8698 => "11111111",
		8699 => "11111111",
		8700 => "11111111",
		8701 => "11111111",
		8702 => "11111111",
		8703 => "11111111",
		8704 => "11111111",
		8705 => "11111111",
		8706 => "11111111",
		8707 => "11111001",
		8708 => "01010011",
		8709 => "11110011",
		8710 => "11111111",
		8711 => "11101110",
		8712 => "01011001",
		8713 => "01000111",
		8714 => "10100011",
		8715 => "11111111",
		8716 => "11111111",
		8717 => "11111111",
		8718 => "10111010",
		8719 => "10100011",
		8720 => "11111111",
		8721 => "11111111",
		8722 => "11111111",
		8723 => "11111111",
		8724 => "11111111",
		8725 => "11111111",
		8726 => "11111111",
		8727 => "11111111",
		8728 => "01101010",
		8729 => "01111100",
		8730 => "11111111",
		8731 => "11111111",
		8732 => "11111111",
		8733 => "11111111",
		8734 => "11111111",
		8735 => "01101010",
		8736 => "01111100",
		8737 => "11111111",
		8738 => "11111111",
		8739 => "11111111",
		8740 => "11110011",
		8741 => "01000111",
		8742 => "10011110",
		8743 => "11111111",
		8744 => "11111111",
		8745 => "11010111",
		8746 => "01000111",
		8747 => "11000101",
		8748 => "11111111",
		8749 => "11111111",
		8750 => "11111111",
		8751 => "11001011",
		8752 => "10100011",
		8753 => "11101000",
		8754 => "11101000",
		8755 => "01000111",
		8756 => "10101110",
		8757 => "11111111",
		8758 => "11111111",
		8759 => "11111111",
		8760 => "11111111",
		8761 => "11111111",
		8762 => "11111111",
		8763 => "11111111",
		8764 => "11111111",
		8765 => "10100011",
		8766 => "11101000",
		8767 => "11111111",
		8768 => "11111111",
		8769 => "11111111",
		8770 => "11111111",
		8771 => "11111111",
		8772 => "11111111",
		8773 => "11111111",
		8774 => "11111111",
		8775 => "11111111",
		8776 => "11111111",
		8777 => "11111111",
		8778 => "11111111",
		8779 => "11111111",
		8780 => "11101110",
		8781 => "01000111",
		8782 => "10100011",
		8783 => "10110100",
		8784 => "10001100",
		8785 => "11101000",
		8786 => "11111111",
		8787 => "11111111",
		8788 => "11111111",
		8789 => "11001011",
		8790 => "01000111",
		8791 => "11000101",
		8792 => "11111111",
		8793 => "11111111",
		8794 => "10101110",
		8795 => "01000111",
		8796 => "11101000",
		8797 => "11111111",
		8798 => "11111111",
		8799 => "11111111",
		8800 => "10010011",
		8801 => "01001101",
		8802 => "11111111",
		8803 => "11111111",
		8804 => "11111111",
		8805 => "11111111",
		8806 => "11111111",
		8807 => "10000111",
		8808 => "01011110",
		8809 => "11111111",
		8810 => "11111111",
		8811 => "11111111",
		8812 => "11111111",
		8813 => "11111111",
		8814 => "11111111",
		8815 => "11111111",
		8816 => "11111111",
		8817 => "11010001",
		8818 => "10011000",
		8819 => "11111111",
		8820 => "11111111",
		8821 => "11111111",
		8822 => "11111111",
		8823 => "11111111",
		8824 => "11111111",
		8825 => "11111111",
		8826 => "11111111",
		8827 => "11111111",
		8828 => "11111111",
		8829 => "11111111",
		8830 => "11111111",
		8831 => "11111111",
		8832 => "11111111",
		8833 => "11111111",
		8834 => "11111111",
		8835 => "11111111",
		8836 => "10010011",
		8837 => "01001101",
		8838 => "10000111",
		8839 => "01011110",
		8840 => "01000111",
		8841 => "01110000",
		8842 => "11111001",
		8843 => "11111111",
		8844 => "11111111",
		8845 => "11000000",
		8846 => "01110000",
		8847 => "11000000",
		8848 => "11111111",
		8849 => "11111111",
		8850 => "11111111",
		8851 => "11111111",
		8852 => "11111111",
		8853 => "11111111",
		8854 => "11111111",
		8855 => "11111111",
		8856 => "01111100",
		8857 => "01101010",
		8858 => "11111111",
		8859 => "11111111",
		8860 => "11111111",
		8861 => "11111111",
		8862 => "11111111",
		8863 => "10001100",
		8864 => "01010011",
		8865 => "11111111",
		8866 => "11111111",
		8867 => "11111111",
		8868 => "11111111",
		8869 => "01101010",
		8870 => "01110000",
		8871 => "10110100",
		8872 => "01111100",
		8873 => "01110000",
		8874 => "01000111",
		8875 => "01100100",
		8876 => "10011110",
		8877 => "11010111",
		8878 => "11111111",
		8879 => "11111111",
		8880 => "11111111",
		8881 => "11111111",
		8882 => "11111001",
		8883 => "01000111",
		8884 => "10100011",
		8885 => "11111111",
		8886 => "11111111",
		8887 => "11111111",
		8888 => "11111111",
		8889 => "11111111",
		8890 => "11111111",
		8891 => "11111111",
		8892 => "11111111",
		8893 => "10011110",
		8894 => "10010011",
		8895 => "01110101",
		8896 => "10100011",
		8897 => "10011000",
		8898 => "10011000",
		8899 => "11101000",
		8900 => "11111111",
		8901 => "11111111",
		8902 => "11111111",
		8903 => "11111111",
		8904 => "11111111",
		8905 => "11111111",
		8906 => "11111111",
		8907 => "11111111",
		8908 => "11000101",
		8909 => "01000111",
		8910 => "11010111",
		8911 => "11111111",
		8912 => "11111111",
		8913 => "11111111",
		8914 => "11111111",
		8915 => "11101110",
		8916 => "10110100",
		8917 => "01110101",
		8918 => "01000111",
		8919 => "01110000",
		8920 => "10100011",
		8921 => "11011100",
		8922 => "10000111",
		8923 => "01010011",
		8924 => "11111111",
		8925 => "11111111",
		8926 => "11111111",
		8927 => "11111111",
		8928 => "01101010",
		8929 => "01110101",
		8930 => "11111111",
		8931 => "11111111",
		8932 => "11111111",
		8933 => "11111111",
		8934 => "11111111",
		8935 => "01110101",
		8936 => "01110101",
		8937 => "11111111",
		8938 => "11111111",
		8939 => "11111111",
		8940 => "11111111",
		8941 => "11111111",
		8942 => "11111111",
		8943 => "11111111",
		8944 => "11111111",
		8945 => "11111111",
		8946 => "11111111",
		8947 => "11111111",
		8948 => "11111111",
		8949 => "11111111",
		8950 => "11111111",
		8951 => "11111111",
		8952 => "11111111",
		8953 => "11111111",
		8954 => "11111111",
		8955 => "11111111",
		8956 => "11111111",
		8957 => "11111111",
		8958 => "11111111",
		8959 => "11111111",
		8960 => "11111111",
		8961 => "11111111",
		8962 => "11111111",
		8963 => "11111111",
		8964 => "11111001",
		8965 => "10011110",
		8966 => "01101010",
		8967 => "01011110",
		8968 => "10010011",
		8969 => "11110011",
		8970 => "11111111",
		8971 => "11111111",
		8972 => "11111111",
		8973 => "01110101",
		8974 => "01110101",
		8975 => "11100010",
		8976 => "11111111",
		8977 => "11111111",
		8978 => "11111111",
		8979 => "11111111",
		8980 => "11111111",
		8981 => "11111111",
		8982 => "11111111",
		8983 => "11111111",
		8984 => "10001100",
		8985 => "01011001",
		8986 => "11111111",
		8987 => "11111111",
		8988 => "11111111",
		8989 => "11111111",
		8990 => "11111111",
		8991 => "10101110",
		8992 => "01000111",
		8993 => "11111111",
		8994 => "11111111",
		8995 => "11111111",
		8996 => "11111111",
		8997 => "10001100",
		8998 => "01000111",
		8999 => "01000111",
		9000 => "01100100",
		9001 => "01110101",
		9002 => "01110101",
		9003 => "01110101",
		9004 => "01001101",
		9005 => "01000111",
		9006 => "10000001",
		9007 => "11101110",
		9008 => "11111111",
		9009 => "11111111",
		9010 => "11111111",
		9011 => "01001101",
		9012 => "10100011",
		9013 => "11111111",
		9014 => "11111111",
		9015 => "11111111",
		9016 => "11111111",
		9017 => "11111111",
		9018 => "11111111",
		9019 => "11111111",
		9020 => "11111111",
		9021 => "11101000",
		9022 => "01101010",
		9023 => "01011110",
		9024 => "01000111",
		9025 => "01000111",
		9026 => "01011001",
		9027 => "10010011",
		9028 => "11111111",
		9029 => "11111111",
		9030 => "11111111",
		9031 => "11111111",
		9032 => "11111111",
		9033 => "11111111",
		9034 => "11111111",
		9035 => "11111111",
		9036 => "10100011",
		9037 => "01000111",
		9038 => "11111001",
		9039 => "11111111",
		9040 => "11111111",
		9041 => "11111001",
		9042 => "10011000",
		9043 => "01001101",
		9044 => "01000111",
		9045 => "01011001",
		9046 => "01110101",
		9047 => "01110000",
		9048 => "01000111",
		9049 => "01000111",
		9050 => "01001101",
		9051 => "10000001",
		9052 => "11111111",
		9053 => "11111111",
		9054 => "11111111",
		9055 => "11110011",
		9056 => "01000111",
		9057 => "10011000",
		9058 => "11111111",
		9059 => "11111111",
		9060 => "11111111",
		9061 => "11111111",
		9062 => "11111111",
		9063 => "01100100",
		9064 => "10000001",
		9065 => "11111111",
		9066 => "11111111",
		9067 => "11111111",
		9068 => "11111111",
		9069 => "11111111",
		9070 => "11111111",
		9071 => "11111111",
		9072 => "11111111",
		9073 => "11111111",
		9074 => "11111111",
		9075 => "11111111",
		9076 => "11111111",
		9077 => "11111111",
		9078 => "11111111",
		9079 => "11111111",
		9080 => "11111111",
		9081 => "11111111",
		9082 => "10101001",
		9083 => "11000101",
		9084 => "11011100",
		9085 => "11111111",
		9086 => "11111111",
		9087 => "11111111",
		9088 => "11111111",
		9089 => "11111111",
		9090 => "11111111",
		9091 => "11111111",
		9092 => "11111111",
		9093 => "11111111",
		9094 => "11111111",
		9095 => "11111111",
		9096 => "11111111",
		9097 => "11111111",
		9098 => "11111111",
		9099 => "11111111",
		9100 => "11111111",
		9101 => "11111111",
		9102 => "11111111",
		9103 => "11111111",
		9104 => "11111111",
		9105 => "11111111",
		9106 => "11111111",
		9107 => "11111111",
		9108 => "11111111",
		9109 => "11111111",
		9110 => "11111111",
		9111 => "11111111",
		9112 => "10101110",
		9113 => "01000111",
		9114 => "11101110",
		9115 => "11111111",
		9116 => "11111111",
		9117 => "11111111",
		9118 => "11111111",
		9119 => "11010111",
		9120 => "01000111",
		9121 => "11111111",
		9122 => "11111111",
		9123 => "11111111",
		9124 => "11111111",
		9125 => "01110000",
		9126 => "01010011",
		9127 => "11001011",
		9128 => "11111111",
		9129 => "11111111",
		9130 => "11111111",
		9131 => "11111111",
		9132 => "11101110",
		9133 => "10100011",
		9134 => "01001101",
		9135 => "01011110",
		9136 => "11101000",
		9137 => "11111111",
		9138 => "11111111",
		9139 => "01100100",
		9140 => "01110101",
		9141 => "11111111",
		9142 => "11111111",
		9143 => "11111111",
		9144 => "11111111",
		9145 => "11111111",
		9146 => "11111111",
		9147 => "11111111",
		9148 => "11111111",
		9149 => "11111111",
		9150 => "11111111",
		9151 => "11111111",
		9152 => "11011100",
		9153 => "11110011",
		9154 => "11111111",
		9155 => "11111111",
		9156 => "11111111",
		9157 => "11111111",
		9158 => "11111111",
		9159 => "11111111",
		9160 => "11111111",
		9161 => "11111111",
		9162 => "11111111",
		9163 => "11111111",
		9164 => "01111100",
		9165 => "01101010",
		9166 => "11111111",
		9167 => "11111111",
		9168 => "11110011",
		9169 => "01101010",
		9170 => "01000111",
		9171 => "10001100",
		9172 => "11100010",
		9173 => "11111111",
		9174 => "11111111",
		9175 => "11111111",
		9176 => "11110011",
		9177 => "01111100",
		9178 => "01000111",
		9179 => "10011000",
		9180 => "11111111",
		9181 => "11111111",
		9182 => "11111111",
		9183 => "11010001",
		9184 => "01000111",
		9185 => "11000101",
		9186 => "11111111",
		9187 => "11111111",
		9188 => "11111111",
		9189 => "11111111",
		9190 => "11111001",
		9191 => "01000111",
		9192 => "10011110",
		9193 => "11111111",
		9194 => "11111111",
		9195 => "11111111",
		9196 => "11111111",
		9197 => "11111111",
		9198 => "11111111",
		9199 => "11111111",
		9200 => "11111111",
		9201 => "10110100",
		9202 => "11111111",
		9203 => "11111111",
		9204 => "11111111",
		9205 => "11111111",
		9206 => "11111111",
		9207 => "11111111",
		9208 => "11111111",
		9209 => "11111111",
		9210 => "10110100",
		9211 => "01011001",
		9212 => "01000111",
		9213 => "11111111",
		9214 => "11111111",
		9215 => "11111111",
		9216 => "11111111",
		9217 => "11111111",
		9218 => "11111111",
		9219 => "11111111",
		9220 => "11111111",
		9221 => "11111111",
		9222 => "11111111",
		9223 => "11111111",
		9224 => "11111111",
		9225 => "11111111",
		9226 => "11111111",
		9227 => "11111111",
		9228 => "11111111",
		9229 => "11111111",
		9230 => "11111111",
		9231 => "11111111",
		9232 => "11111111",
		9233 => "11111111",
		9234 => "11111111",
		9235 => "11111111",
		9236 => "11111111",
		9237 => "11111111",
		9238 => "11111111",
		9239 => "11111111",
		9240 => "11010001",
		9241 => "01000111",
		9242 => "11000101",
		9243 => "11111111",
		9244 => "11111111",
		9245 => "11111111",
		9246 => "11111111",
		9247 => "11111001",
		9248 => "01001101",
		9249 => "11111111",
		9250 => "11111111",
		9251 => "11111111",
		9252 => "11000000",
		9253 => "01000111",
		9254 => "10110100",
		9255 => "11111111",
		9256 => "11111111",
		9257 => "11111111",
		9258 => "11111111",
		9259 => "11111111",
		9260 => "11111111",
		9261 => "11111111",
		9262 => "11010001",
		9263 => "01010011",
		9264 => "01101010",
		9265 => "11111111",
		9266 => "11111111",
		9267 => "10100011",
		9268 => "01000111",
		9269 => "11101000",
		9270 => "11111111",
		9271 => "11111111",
		9272 => "11111111",
		9273 => "11111111",
		9274 => "11111111",
		9275 => "11111111",
		9276 => "11111111",
		9277 => "11111111",
		9278 => "11111111",
		9279 => "11111111",
		9280 => "11111111",
		9281 => "11111111",
		9282 => "11111111",
		9283 => "11111111",
		9284 => "11111111",
		9285 => "11111111",
		9286 => "11111111",
		9287 => "11111111",
		9288 => "11111111",
		9289 => "11111111",
		9290 => "11111111",
		9291 => "11100010",
		9292 => "01000111",
		9293 => "10100011",
		9294 => "11111111",
		9295 => "11111001",
		9296 => "01110000",
		9297 => "01000111",
		9298 => "11001011",
		9299 => "11111111",
		9300 => "11111111",
		9301 => "11111111",
		9302 => "11111111",
		9303 => "11111111",
		9304 => "11111111",
		9305 => "11111111",
		9306 => "01110101",
		9307 => "01001101",
		9308 => "11101110",
		9309 => "11111111",
		9310 => "11111111",
		9311 => "10101001",
		9312 => "01000111",
		9313 => "11101110",
		9314 => "11111111",
		9315 => "11111111",
		9316 => "11111111",
		9317 => "11111111",
		9318 => "11010001",
		9319 => "01000111",
		9320 => "11000101",
		9321 => "11111111",
		9322 => "11111111",
		9323 => "11111111",
		9324 => "11111111",
		9325 => "11111111",
		9326 => "11111111",
		9327 => "11111111",
		9328 => "11111111",
		9329 => "01100100",
		9330 => "11111111",
		9331 => "11111111",
		9332 => "11111111",
		9333 => "11111111",
		9334 => "11111111",
		9335 => "11111111",
		9336 => "11111111",
		9337 => "11111111",
		9338 => "11111111",
		9339 => "11110011",
		9340 => "01011110",
		9341 => "11111111",
		9342 => "11111111",
		9343 => "11111111",
		9344 => "11111111",
		9345 => "11111111",
		9346 => "11111111",
		9347 => "11111111",
		9348 => "11111111",
		9349 => "11111111",
		9350 => "11111111",
		9351 => "11111111",
		9352 => "11111111",
		9353 => "11111111",
		9354 => "11111111",
		9355 => "11111111",
		9356 => "11111111",
		9357 => "11111111",
		9358 => "11111111",
		9359 => "11111111",
		9360 => "11111111",
		9361 => "11111111",
		9362 => "11111111",
		9363 => "11111111",
		9364 => "11111111",
		9365 => "11111111",
		9366 => "11111111",
		9367 => "11111111",
		9368 => "11111001",
		9369 => "01000111",
		9370 => "10100011",
		9371 => "11111111",
		9372 => "11111111",
		9373 => "11111111",
		9374 => "11111111",
		9375 => "11111111",
		9376 => "01101010",
		9377 => "11111111",
		9378 => "11111111",
		9379 => "11111111",
		9380 => "01110101",
		9381 => "01101010",
		9382 => "11111111",
		9383 => "11111111",
		9384 => "11111111",
		9385 => "11111111",
		9386 => "11111111",
		9387 => "11111111",
		9388 => "11111111",
		9389 => "11111111",
		9390 => "11111111",
		9391 => "10111010",
		9392 => "01000111",
		9393 => "10101110",
		9394 => "11111111",
		9395 => "11101000",
		9396 => "01000111",
		9397 => "10100011",
		9398 => "11111111",
		9399 => "11111111",
		9400 => "11111111",
		9401 => "11111111",
		9402 => "11111111",
		9403 => "11111111",
		9404 => "11101000",
		9405 => "11111111",
		9406 => "11111111",
		9407 => "10111010",
		9408 => "10100011",
		9409 => "10100011",
		9410 => "11000101",
		9411 => "11111111",
		9412 => "11110011",
		9413 => "11111111",
		9414 => "11111111",
		9415 => "11111111",
		9416 => "11111111",
		9417 => "11111111",
		9418 => "11111111",
		9419 => "10011000",
		9420 => "01001101",
		9421 => "11101110",
		9422 => "11111111",
		9423 => "10010011",
		9424 => "01000111",
		9425 => "10101110",
		9426 => "11111111",
		9427 => "11111111",
		9428 => "11111111",
		9429 => "11111111",
		9430 => "11111111",
		9431 => "11111111",
		9432 => "11111111",
		9433 => "11111111",
		9434 => "11011100",
		9435 => "01000111",
		9436 => "10011000",
		9437 => "11111111",
		9438 => "11111111",
		9439 => "01111100",
		9440 => "01011110",
		9441 => "11111111",
		9442 => "11111111",
		9443 => "11111111",
		9444 => "11111111",
		9445 => "11111111",
		9446 => "10101110",
		9447 => "01000111",
		9448 => "11101000",
		9449 => "11111111",
		9450 => "11111111",
		9451 => "11111111",
		9452 => "11111111",
		9453 => "11111111",
		9454 => "11111111",
		9455 => "11111111",
		9456 => "11110011",
		9457 => "01000111",
		9458 => "10011000",
		9459 => "11010001",
		9460 => "11110011",
		9461 => "11111111",
		9462 => "11111111",
		9463 => "11111111",
		9464 => "11111111",
		9465 => "11111111",
		9466 => "11111111",
		9467 => "11101110",
		9468 => "01110000",
		9469 => "11111111",
		9470 => "11111111",
		9471 => "11111111",
		9472 => "11111111",
		9473 => "11111111",
		9474 => "11111111",
		9475 => "11111111",
		9476 => "11111111",
		9477 => "11111111",
		9478 => "11111111",
		9479 => "11111111",
		9480 => "11111111",
		9481 => "11111111",
		9482 => "11111111",
		9483 => "11111111",
		9484 => "11111111",
		9485 => "11111111",
		9486 => "11111111",
		9487 => "11111111",
		9488 => "11111111",
		9489 => "11111111",
		9490 => "11111111",
		9491 => "11111111",
		9492 => "11111111",
		9493 => "11111111",
		9494 => "11111111",
		9495 => "11111111",
		9496 => "11111111",
		9497 => "10010011",
		9498 => "01010011",
		9499 => "11111111",
		9500 => "11111111",
		9501 => "11111111",
		9502 => "11111111",
		9503 => "11111111",
		9504 => "11101000",
		9505 => "10101110",
		9506 => "11111111",
		9507 => "10110100",
		9508 => "01001101",
		9509 => "11110011",
		9510 => "11111111",
		9511 => "11111111",
		9512 => "11111111",
		9513 => "11111111",
		9514 => "11111111",
		9515 => "11111111",
		9516 => "11111111",
		9517 => "11111111",
		9518 => "11111111",
		9519 => "11111111",
		9520 => "11101110",
		9521 => "01011001",
		9522 => "01011110",
		9523 => "11101110",
		9524 => "11000101",
		9525 => "01000111",
		9526 => "11111111",
		9527 => "11111111",
		9528 => "11111111",
		9529 => "11111111",
		9530 => "11111001",
		9531 => "11010001",
		9532 => "10110100",
		9533 => "01110101",
		9534 => "01111100",
		9535 => "10011110",
		9536 => "01110101",
		9537 => "10011110",
		9538 => "01111100",
		9539 => "01111100",
		9540 => "10101001",
		9541 => "10100011",
		9542 => "11101000",
		9543 => "11111111",
		9544 => "11111111",
		9545 => "11111111",
		9546 => "10011000",
		9547 => "01000111",
		9548 => "11011100",
		9549 => "11101000",
		9550 => "01010011",
		9551 => "01110000",
		9552 => "11111001",
		9553 => "11111111",
		9554 => "11111111",
		9555 => "11111111",
		9556 => "11111111",
		9557 => "11111111",
		9558 => "11111111",
		9559 => "11111111",
		9560 => "11111111",
		9561 => "11111111",
		9562 => "11111111",
		9563 => "10111010",
		9564 => "01000111",
		9565 => "11011100",
		9566 => "10111010",
		9567 => "01000111",
		9568 => "11010001",
		9569 => "11111111",
		9570 => "11111111",
		9571 => "11111111",
		9572 => "11111111",
		9573 => "11111111",
		9574 => "01011110",
		9575 => "10000001",
		9576 => "11111111",
		9577 => "11111111",
		9578 => "11111111",
		9579 => "11111111",
		9580 => "11111111",
		9581 => "11111111",
		9582 => "11111111",
		9583 => "11111111",
		9584 => "10110100",
		9585 => "10001100",
		9586 => "11010001",
		9587 => "10011110",
		9588 => "01110101",
		9589 => "01011110",
		9590 => "01000111",
		9591 => "01000111",
		9592 => "01000111",
		9593 => "01000111",
		9594 => "01000111",
		9595 => "01000111",
		9596 => "10101110",
		9597 => "11111111",
		9598 => "11111111",
		9599 => "11111111",
		9600 => "11111111",
		9601 => "11111111",
		9602 => "11111111",
		9603 => "11111111",
		9604 => "11111111",
		9605 => "11111111",
		9606 => "11111111",
		9607 => "11111111",
		9608 => "11111111",
		9609 => "11111111",
		9610 => "11111111",
		9611 => "11111111",
		9612 => "11111111",
		9613 => "11111111",
		9614 => "11111111",
		9615 => "11111111",
		9616 => "11111111",
		9617 => "11111111",
		9618 => "11111111",
		9619 => "11111111",
		9620 => "11111111",
		9621 => "11111111",
		9622 => "11111111",
		9623 => "11111111",
		9624 => "11111111",
		9625 => "11000000",
		9626 => "01000111",
		9627 => "11010001",
		9628 => "11111111",
		9629 => "11111111",
		9630 => "11111111",
		9631 => "11111111",
		9632 => "11111111",
		9633 => "01101010",
		9634 => "11111111",
		9635 => "10001100",
		9636 => "01011110",
		9637 => "11111111",
		9638 => "11111111",
		9639 => "11111111",
		9640 => "11111111",
		9641 => "11111111",
		9642 => "11111111",
		9643 => "11111111",
		9644 => "11111111",
		9645 => "11111111",
		9646 => "11111111",
		9647 => "11111111",
		9648 => "11111111",
		9649 => "10101110",
		9650 => "01000111",
		9651 => "01001101",
		9652 => "01110101",
		9653 => "01000111",
		9654 => "11110011",
		9655 => "11111111",
		9656 => "11111111",
		9657 => "11111111",
		9658 => "11111111",
		9659 => "11111111",
		9660 => "11111111",
		9661 => "11111111",
		9662 => "11111111",
		9663 => "11111111",
		9664 => "11111111",
		9665 => "11111111",
		9666 => "11111111",
		9667 => "11111111",
		9668 => "11111111",
		9669 => "11111111",
		9670 => "11111111",
		9671 => "11111111",
		9672 => "11111111",
		9673 => "11111111",
		9674 => "01000111",
		9675 => "01011110",
		9676 => "10001100",
		9677 => "01001101",
		9678 => "01000111",
		9679 => "11001011",
		9680 => "11111111",
		9681 => "11111111",
		9682 => "11111111",
		9683 => "11111111",
		9684 => "11111111",
		9685 => "11111111",
		9686 => "11111111",
		9687 => "11111111",
		9688 => "11111111",
		9689 => "11111111",
		9690 => "11111111",
		9691 => "11011100",
		9692 => "01000111",
		9693 => "11000000",
		9694 => "01111100",
		9695 => "01011001",
		9696 => "11111111",
		9697 => "11111111",
		9698 => "11111111",
		9699 => "11111111",
		9700 => "11111111",
		9701 => "11100010",
		9702 => "01000111",
		9703 => "10101001",
		9704 => "11111111",
		9705 => "11111111",
		9706 => "11111111",
		9707 => "11111111",
		9708 => "11111111",
		9709 => "11111111",
		9710 => "11111111",
		9711 => "11111111",
		9712 => "10011110",
		9713 => "11101110",
		9714 => "11111111",
		9715 => "11111111",
		9716 => "11111111",
		9717 => "11111111",
		9718 => "11111111",
		9719 => "11010001",
		9720 => "11000000",
		9721 => "10100011",
		9722 => "01111100",
		9723 => "01010011",
		9724 => "11001011",
		9725 => "11111111",
		9726 => "11111111",
		9727 => "11111111",
		9728 => "11111111",
		9729 => "11111111",
		9730 => "11111111",
		9731 => "11111111",
		9732 => "11111111",
		9733 => "11111111",
		9734 => "11111111",
		9735 => "11111111",
		9736 => "11111111",
		9737 => "11111111",
		9738 => "11111111",
		9739 => "11111111",
		9740 => "11111111",
		9741 => "11111111",
		9742 => "11111111",
		9743 => "11111111",
		9744 => "11111111",
		9745 => "11111111",
		9746 => "11111111",
		9747 => "11111111",
		9748 => "11111111",
		9749 => "11111111",
		9750 => "11111111",
		9751 => "11111111",
		9752 => "11111111",
		9753 => "11111001",
		9754 => "01001101",
		9755 => "10011000",
		9756 => "11111111",
		9757 => "11111111",
		9758 => "11111111",
		9759 => "11111111",
		9760 => "11111111",
		9761 => "01000111",
		9762 => "11011100",
		9763 => "10001100",
		9764 => "01101010",
		9765 => "11111111",
		9766 => "11111111",
		9767 => "11111111",
		9768 => "11111111",
		9769 => "11111111",
		9770 => "11111111",
		9771 => "11111111",
		9772 => "11111111",
		9773 => "11111111",
		9774 => "11111111",
		9775 => "11111111",
		9776 => "11111111",
		9777 => "11011100",
		9778 => "01000111",
		9779 => "01110000",
		9780 => "01110101",
		9781 => "10100011",
		9782 => "01101010",
		9783 => "11110011",
		9784 => "11111111",
		9785 => "11111111",
		9786 => "11111111",
		9787 => "11111111",
		9788 => "11111111",
		9789 => "11111111",
		9790 => "11010111",
		9791 => "01110101",
		9792 => "10100011",
		9793 => "10011000",
		9794 => "10110100",
		9795 => "11111111",
		9796 => "11111111",
		9797 => "11111111",
		9798 => "11111111",
		9799 => "11111111",
		9800 => "11111111",
		9801 => "11001011",
		9802 => "01011110",
		9803 => "01110101",
		9804 => "01011110",
		9805 => "01011001",
		9806 => "01001101",
		9807 => "11111111",
		9808 => "11111111",
		9809 => "11111111",
		9810 => "11111111",
		9811 => "11111111",
		9812 => "11111111",
		9813 => "11111111",
		9814 => "11111111",
		9815 => "11111111",
		9816 => "11111111",
		9817 => "11111111",
		9818 => "11111111",
		9819 => "11101110",
		9820 => "01000111",
		9821 => "10111010",
		9822 => "01001101",
		9823 => "10011000",
		9824 => "11111111",
		9825 => "11111111",
		9826 => "11111111",
		9827 => "11111111",
		9828 => "11111111",
		9829 => "10100011",
		9830 => "01000111",
		9831 => "11101000",
		9832 => "11111111",
		9833 => "11111111",
		9834 => "11111111",
		9835 => "11111111",
		9836 => "11111111",
		9837 => "11111111",
		9838 => "11111111",
		9839 => "11111111",
		9840 => "11111111",
		9841 => "11111111",
		9842 => "11111111",
		9843 => "11111111",
		9844 => "11111111",
		9845 => "11111111",
		9846 => "11111111",
		9847 => "11111111",
		9848 => "11111111",
		9849 => "11111111",
		9850 => "11111111",
		9851 => "01101010",
		9852 => "11101110",
		9853 => "11111111",
		9854 => "11111111",
		9855 => "11111111",
		9856 => "11111111",
		9857 => "11111111",
		9858 => "11111111",
		9859 => "11111111",
		9860 => "11111111",
		9861 => "11111111",
		9862 => "11111111",
		9863 => "11111111",
		9864 => "11111111",
		9865 => "11111111",
		9866 => "11111111",
		9867 => "11111111",
		9868 => "11111111",
		9869 => "11111111",
		9870 => "11111111",
		9871 => "11111111",
		9872 => "11111111",
		9873 => "11111111",
		9874 => "11111111",
		9875 => "11111111",
		9876 => "11111111",
		9877 => "11111111",
		9878 => "11111111",
		9879 => "11111111",
		9880 => "11111111",
		9881 => "11111111",
		9882 => "10000111",
		9883 => "01011110",
		9884 => "11111111",
		9885 => "11111111",
		9886 => "11111111",
		9887 => "11111111",
		9888 => "11111111",
		9889 => "01001101",
		9890 => "10000001",
		9891 => "10001100",
		9892 => "01110000",
		9893 => "11111111",
		9894 => "11111111",
		9895 => "11111111",
		9896 => "11111111",
		9897 => "11111111",
		9898 => "11111111",
		9899 => "11111111",
		9900 => "11111111",
		9901 => "11111111",
		9902 => "11111111",
		9903 => "11111111",
		9904 => "11111111",
		9905 => "11000000",
		9906 => "01000111",
		9907 => "11010001",
		9908 => "11111111",
		9909 => "11111111",
		9910 => "01001101",
		9911 => "01101010",
		9912 => "11100010",
		9913 => "11111111",
		9914 => "11111111",
		9915 => "11111111",
		9916 => "11111111",
		9917 => "11111111",
		9918 => "11111111",
		9919 => "11100010",
		9920 => "10101001",
		9921 => "10011110",
		9922 => "10111010",
		9923 => "11111111",
		9924 => "11111111",
		9925 => "11111111",
		9926 => "11111111",
		9927 => "11111111",
		9928 => "11000000",
		9929 => "01001101",
		9930 => "11110011",
		9931 => "11111111",
		9932 => "11111111",
		9933 => "10100011",
		9934 => "01001101",
		9935 => "11101110",
		9936 => "11111111",
		9937 => "11111111",
		9938 => "11111111",
		9939 => "11111111",
		9940 => "11111111",
		9941 => "11111111",
		9942 => "11111111",
		9943 => "11111111",
		9944 => "11111111",
		9945 => "11111111",
		9946 => "11111111",
		9947 => "11111001",
		9948 => "01000111",
		9949 => "10111010",
		9950 => "01000111",
		9951 => "11011100",
		9952 => "11111111",
		9953 => "11111111",
		9954 => "11111111",
		9955 => "11111111",
		9956 => "11111111",
		9957 => "01100100",
		9958 => "01100100",
		9959 => "11111111",
		9960 => "11111111",
		9961 => "11111111",
		9962 => "11111111",
		9963 => "11111111",
		9964 => "11111111",
		9965 => "11111111",
		9966 => "11111111",
		9967 => "11111111",
		9968 => "11111111",
		9969 => "11111111",
		9970 => "11111111",
		9971 => "11111111",
		9972 => "11111111",
		9973 => "11111111",
		9974 => "11111111",
		9975 => "11111111",
		9976 => "11111111",
		9977 => "11111111",
		9978 => "11111111",
		9979 => "01011001",
		9980 => "11111111",
		9981 => "11111111",
		9982 => "11111111",
		9983 => "11111111",
		9984 => "11111111",
		9985 => "11111111",
		9986 => "11111111",
		9987 => "11111111",
		9988 => "11111111",
		9989 => "11111111",
		9990 => "11111111",
		9991 => "11111111",
		9992 => "11111111",
		9993 => "11111111",
		9994 => "11111111",
		9995 => "11111111",
		9996 => "11111111",
		9997 => "11111111",
		9998 => "11111111",
		9999 => "11111111",
		10000 => "11111111",
		10001 => "11101110",
		10002 => "11111111",
		10003 => "11111111",
		10004 => "11111111",
		10005 => "11111111",
		10006 => "11111111",
		10007 => "11111111",
		10008 => "11111111",
		10009 => "11111111",
		10010 => "11000000",
		10011 => "01000111",
		10012 => "11010111",
		10013 => "11111111",
		10014 => "11111111",
		10015 => "11111111",
		10016 => "11111111",
		10017 => "10011000",
		10018 => "01001101",
		10019 => "10010011",
		10020 => "01010011",
		10021 => "11111111",
		10022 => "11111111",
		10023 => "11111111",
		10024 => "11111111",
		10025 => "11111111",
		10026 => "11111111",
		10027 => "11111111",
		10028 => "11111111",
		10029 => "11111111",
		10030 => "11111111",
		10031 => "11111111",
		10032 => "11010111",
		10033 => "01100100",
		10034 => "01011001",
		10035 => "11111001",
		10036 => "11110011",
		10037 => "01111100",
		10038 => "11010001",
		10039 => "01011001",
		10040 => "01010011",
		10041 => "10011110",
		10042 => "11101000",
		10043 => "11111111",
		10044 => "11111111",
		10045 => "11111111",
		10046 => "11111111",
		10047 => "11111111",
		10048 => "11111111",
		10049 => "11111111",
		10050 => "11111111",
		10051 => "11111111",
		10052 => "11111111",
		10053 => "11111111",
		10054 => "11110011",
		10055 => "10001100",
		10056 => "01000111",
		10057 => "01110000",
		10058 => "11010001",
		10059 => "10100011",
		10060 => "11111111",
		10061 => "11010001",
		10062 => "01000111",
		10063 => "10011110",
		10064 => "11111001",
		10065 => "11111111",
		10066 => "11111111",
		10067 => "11111111",
		10068 => "11111111",
		10069 => "11111111",
		10070 => "11111111",
		10071 => "11111111",
		10072 => "11111111",
		10073 => "11111111",
		10074 => "11111111",
		10075 => "11011100",
		10076 => "01000111",
		10077 => "11000000",
		10078 => "01101010",
		10079 => "11111111",
		10080 => "11111111",
		10081 => "11111111",
		10082 => "11111111",
		10083 => "11111111",
		10084 => "11100010",
		10085 => "01000111",
		10086 => "10100011",
		10087 => "11111111",
		10088 => "11111111",
		10089 => "11111111",
		10090 => "11111111",
		10091 => "11111111",
		10092 => "11111111",
		10093 => "11111111",
		10094 => "11111111",
		10095 => "11111111",
		10096 => "11111111",
		10097 => "11111111",
		10098 => "11111111",
		10099 => "11111111",
		10100 => "11111111",
		10101 => "11111111",
		10102 => "11111111",
		10103 => "11111111",
		10104 => "11111111",
		10105 => "11010111",
		10106 => "10100011",
		10107 => "01110000",
		10108 => "11111111",
		10109 => "11111111",
		10110 => "11111111",
		10111 => "11111111",
		10112 => "11111111",
		10113 => "11111111",
		10114 => "11111111",
		10115 => "11111111",
		10116 => "11111111",
		10117 => "11111111",
		10118 => "11111111",
		10119 => "11111111",
		10120 => "11111111",
		10121 => "11111111",
		10122 => "11111111",
		10123 => "11111111",
		10124 => "11111111",
		10125 => "11111111",
		10126 => "11101000",
		10127 => "10100011",
		10128 => "01011110",
		10129 => "10011110",
		10130 => "11111111",
		10131 => "11111111",
		10132 => "11111111",
		10133 => "11111111",
		10134 => "11111111",
		10135 => "11111111",
		10136 => "11111111",
		10137 => "11111111",
		10138 => "11111001",
		10139 => "01001101",
		10140 => "10011000",
		10141 => "11111111",
		10142 => "11111111",
		10143 => "11111111",
		10144 => "11111111",
		10145 => "11101110",
		10146 => "01001101",
		10147 => "01001101",
		10148 => "01000111",
		10149 => "11101110",
		10150 => "11111111",
		10151 => "11111111",
		10152 => "11111111",
		10153 => "11111111",
		10154 => "11111111",
		10155 => "11111111",
		10156 => "11111111",
		10157 => "11111111",
		10158 => "10001100",
		10159 => "01000111",
		10160 => "01000111",
		10161 => "01010011",
		10162 => "11010001",
		10163 => "11111111",
		10164 => "11111001",
		10165 => "01011110",
		10166 => "11110011",
		10167 => "11110011",
		10168 => "10010011",
		10169 => "01000111",
		10170 => "01000111",
		10171 => "10000001",
		10172 => "11011100",
		10173 => "11111111",
		10174 => "11111111",
		10175 => "11111111",
		10176 => "11111111",
		10177 => "11111111",
		10178 => "11111111",
		10179 => "11111111",
		10180 => "11111111",
		10181 => "11001011",
		10182 => "01011001",
		10183 => "01000111",
		10184 => "10011110",
		10185 => "11111001",
		10186 => "01001101",
		10187 => "01111100",
		10188 => "11111111",
		10189 => "11111111",
		10190 => "10010011",
		10191 => "01000111",
		10192 => "01010011",
		10193 => "01110101",
		10194 => "11001011",
		10195 => "11111111",
		10196 => "11111111",
		10197 => "11111111",
		10198 => "11111111",
		10199 => "11111111",
		10200 => "11111111",
		10201 => "11111111",
		10202 => "11111111",
		10203 => "11000000",
		10204 => "01000111",
		10205 => "10101001",
		10206 => "10110100",
		10207 => "11111111",
		10208 => "11111111",
		10209 => "11111111",
		10210 => "11111111",
		10211 => "11111111",
		10212 => "10100011",
		10213 => "01000111",
		10214 => "11100010",
		10215 => "11111111",
		10216 => "11111111",
		10217 => "11111111",
		10218 => "11111111",
		10219 => "11111111",
		10220 => "11111111",
		10221 => "11111111",
		10222 => "11111111",
		10223 => "10100011",
		10224 => "11111111",
		10225 => "11111111",
		10226 => "11111111",
		10227 => "11111111",
		10228 => "11111111",
		10229 => "11111111",
		10230 => "11111111",
		10231 => "11111111",
		10232 => "10110100",
		10233 => "01110101",
		10234 => "01000111",
		10235 => "10010011",
		10236 => "11111111",
		10237 => "11111111",
		10238 => "11111111",
		10239 => "11111111",
		10240 => "11111111",
		10241 => "11111111",
		10242 => "11111111",
		10243 => "11111111",
		10244 => "11111111",
		10245 => "11111111",
		10246 => "11111111",
		10247 => "11111111",
		10248 => "11111111",
		10249 => "11111111",
		10250 => "11111111",
		10251 => "11111111",
		10252 => "11111001",
		10253 => "01111100",
		10254 => "01000111",
		10255 => "01000111",
		10256 => "01011110",
		10257 => "11111001",
		10258 => "11111111",
		10259 => "11111111",
		10260 => "11111111",
		10261 => "11111111",
		10262 => "11111111",
		10263 => "11111111",
		10264 => "11111111",
		10265 => "11111111",
		10266 => "11111111",
		10267 => "10011000",
		10268 => "01001101",
		10269 => "11101110",
		10270 => "11111111",
		10271 => "11111111",
		10272 => "11111111",
		10273 => "11111111",
		10274 => "10010011",
		10275 => "01000111",
		10276 => "01000111",
		10277 => "11000000",
		10278 => "11111111",
		10279 => "11111111",
		10280 => "11111111",
		10281 => "11111111",
		10282 => "11111111",
		10283 => "11111111",
		10284 => "11111111",
		10285 => "11111111",
		10286 => "01100100",
		10287 => "01100100",
		10288 => "10101001",
		10289 => "11101000",
		10290 => "11111111",
		10291 => "11111111",
		10292 => "11111111",
		10293 => "11001011",
		10294 => "11000101",
		10295 => "11111111",
		10296 => "11111111",
		10297 => "11101000",
		10298 => "10011000",
		10299 => "01010011",
		10300 => "01000111",
		10301 => "10000001",
		10302 => "11011100",
		10303 => "11011100",
		10304 => "11000000",
		10305 => "11010001",
		10306 => "10110100",
		10307 => "11100010",
		10308 => "01111100",
		10309 => "01000111",
		10310 => "01100100",
		10311 => "11010111",
		10312 => "11111111",
		10313 => "11111111",
		10314 => "01001101",
		10315 => "11110011",
		10316 => "11111111",
		10317 => "11111111",
		10318 => "11111111",
		10319 => "11001011",
		10320 => "10011000",
		10321 => "01001101",
		10322 => "10010011",
		10323 => "11111111",
		10324 => "11111111",
		10325 => "11111111",
		10326 => "11111111",
		10327 => "11111111",
		10328 => "11111111",
		10329 => "11111111",
		10330 => "11111111",
		10331 => "10010011",
		10332 => "01001101",
		10333 => "01101010",
		10334 => "11111001",
		10335 => "11111111",
		10336 => "11111111",
		10337 => "11111111",
		10338 => "11111111",
		10339 => "11111001",
		10340 => "01011001",
		10341 => "01101010",
		10342 => "11111111",
		10343 => "11111111",
		10344 => "11111111",
		10345 => "11111111",
		10346 => "11111111",
		10347 => "11111111",
		10348 => "11111111",
		10349 => "11111111",
		10350 => "11111001",
		10351 => "01001101",
		10352 => "11111111",
		10353 => "11111111",
		10354 => "11111111",
		10355 => "11111111",
		10356 => "11111111",
		10357 => "11111111",
		10358 => "11111111",
		10359 => "11111111",
		10360 => "11111111",
		10361 => "11111111",
		10362 => "11111111",
		10363 => "11111111",
		10364 => "11111111",
		10365 => "11111111",
		10366 => "11111111",
		10367 => "11111111",
		10368 => "11111111",
		10369 => "11111111",
		10370 => "11111111",
		10371 => "11111111",
		10372 => "11111111",
		10373 => "11111111",
		10374 => "11100010",
		10375 => "11111111",
		10376 => "11111111",
		10377 => "11111111",
		10378 => "11010111",
		10379 => "10001100",
		10380 => "01010011",
		10381 => "10111010",
		10382 => "01011110",
		10383 => "01000111",
		10384 => "11001011",
		10385 => "11111111",
		10386 => "11111111",
		10387 => "11111111",
		10388 => "11111111",
		10389 => "11111111",
		10390 => "11111111",
		10391 => "11111111",
		10392 => "11111111",
		10393 => "11111111",
		10394 => "11111111",
		10395 => "11101110",
		10396 => "01000111",
		10397 => "10011110",
		10398 => "11111111",
		10399 => "11111111",
		10400 => "11111111",
		10401 => "11111111",
		10402 => "11101110",
		10403 => "01001101",
		10404 => "01000111",
		10405 => "01111100",
		10406 => "11111111",
		10407 => "11111111",
		10408 => "11111111",
		10409 => "11111111",
		10410 => "11111111",
		10411 => "11111111",
		10412 => "11111111",
		10413 => "10110100",
		10414 => "01000111",
		10415 => "10100011",
		10416 => "11111111",
		10417 => "11111111",
		10418 => "11111111",
		10419 => "11111111",
		10420 => "11111111",
		10421 => "11011100",
		10422 => "10101110",
		10423 => "11111111",
		10424 => "11111111",
		10425 => "11111111",
		10426 => "11111111",
		10427 => "11110011",
		10428 => "10100011",
		10429 => "01010011",
		10430 => "01000111",
		10431 => "01001101",
		10432 => "01001101",
		10433 => "01000111",
		10434 => "01000111",
		10435 => "01000111",
		10436 => "01010011",
		10437 => "10101110",
		10438 => "11111111",
		10439 => "11111111",
		10440 => "11111111",
		10441 => "11111111",
		10442 => "01011110",
		10443 => "11111111",
		10444 => "11111111",
		10445 => "11111111",
		10446 => "11111111",
		10447 => "11111111",
		10448 => "11111111",
		10449 => "10001100",
		10450 => "01001101",
		10451 => "11011100",
		10452 => "11111111",
		10453 => "11111111",
		10454 => "11111111",
		10455 => "11111111",
		10456 => "11111111",
		10457 => "11111111",
		10458 => "11111001",
		10459 => "01011001",
		10460 => "01000111",
		10461 => "01000111",
		10462 => "11111111",
		10463 => "11111111",
		10464 => "11111111",
		10465 => "11111111",
		10466 => "11111111",
		10467 => "10101110",
		10468 => "01000111",
		10469 => "11000101",
		10470 => "11111111",
		10471 => "11111111",
		10472 => "11111111",
		10473 => "11111111",
		10474 => "11111111",
		10475 => "11111111",
		10476 => "11111111",
		10477 => "11111111",
		10478 => "11000000",
		10479 => "01000111",
		10480 => "01011001",
		10481 => "10010011",
		10482 => "11010001",
		10483 => "11111111",
		10484 => "11111111",
		10485 => "11111111",
		10486 => "11111111",
		10487 => "11111111",
		10488 => "11111111",
		10489 => "11111111",
		10490 => "11111111",
		10491 => "11111111",
		10492 => "11111111",
		10493 => "11111111",
		10494 => "11111111",
		10495 => "11111111",
		10496 => "11111111",
		10497 => "11111111",
		10498 => "11111111",
		10499 => "11111111",
		10500 => "11111111",
		10501 => "11111111",
		10502 => "01110000",
		10503 => "10111010",
		10504 => "10101001",
		10505 => "01011110",
		10506 => "01100100",
		10507 => "10101001",
		10508 => "11101110",
		10509 => "10100011",
		10510 => "01000111",
		10511 => "10001100",
		10512 => "11111111",
		10513 => "11111111",
		10514 => "11111111",
		10515 => "11111111",
		10516 => "11111111",
		10517 => "11111111",
		10518 => "11111111",
		10519 => "11111111",
		10520 => "11111111",
		10521 => "11111111",
		10522 => "11111111",
		10523 => "11111111",
		10524 => "10000001",
		10525 => "01011001",
		10526 => "11111001",
		10527 => "11111111",
		10528 => "11111111",
		10529 => "11111111",
		10530 => "11111111",
		10531 => "10101110",
		10532 => "01000111",
		10533 => "01000111",
		10534 => "11101110",
		10535 => "11111111",
		10536 => "11111111",
		10537 => "11111001",
		10538 => "01011110",
		10539 => "01011110",
		10540 => "01011110",
		10541 => "01000111",
		10542 => "01101010",
		10543 => "11111001",
		10544 => "11111111",
		10545 => "11110011",
		10546 => "11011100",
		10547 => "11111111",
		10548 => "11111001",
		10549 => "10001100",
		10550 => "11010001",
		10551 => "11111111",
		10552 => "11111111",
		10553 => "11111111",
		10554 => "11111111",
		10555 => "11111111",
		10556 => "11111111",
		10557 => "11110011",
		10558 => "01101010",
		10559 => "01000111",
		10560 => "01110101",
		10561 => "01110000",
		10562 => "01000111",
		10563 => "01110000",
		10564 => "11110011",
		10565 => "11111111",
		10566 => "11111111",
		10567 => "11111111",
		10568 => "11111111",
		10569 => "11111111",
		10570 => "01000111",
		10571 => "11010001",
		10572 => "11111111",
		10573 => "11111111",
		10574 => "11111111",
		10575 => "11111111",
		10576 => "11111111",
		10577 => "11101000",
		10578 => "01010011",
		10579 => "01000111",
		10580 => "01101010",
		10581 => "01000111",
		10582 => "10101110",
		10583 => "11111111",
		10584 => "11111111",
		10585 => "11111111",
		10586 => "11000101",
		10587 => "01000111",
		10588 => "01000111",
		10589 => "10000001",
		10590 => "11111111",
		10591 => "11111111",
		10592 => "11111111",
		10593 => "11111111",
		10594 => "11111111",
		10595 => "01011001",
		10596 => "01101010",
		10597 => "11111111",
		10598 => "11111111",
		10599 => "11111111",
		10600 => "11111111",
		10601 => "11111111",
		10602 => "11111111",
		10603 => "11111111",
		10604 => "11111111",
		10605 => "11111111",
		10606 => "10000001",
		10607 => "01101010",
		10608 => "01010011",
		10609 => "01000111",
		10610 => "01000111",
		10611 => "10010011",
		10612 => "11011100",
		10613 => "11111111",
		10614 => "11111111",
		10615 => "11111111",
		10616 => "11111111",
		10617 => "11111111",
		10618 => "11111111",
		10619 => "11111111",
		10620 => "11111111",
		10621 => "11111111",
		10622 => "11111111",
		10623 => "11111111",
		10624 => "11111111",
		10625 => "11111111",
		10626 => "11111111",
		10627 => "11111111",
		10628 => "11111111",
		10629 => "11111111",
		10630 => "10110100",
		10631 => "01001101",
		10632 => "10010011",
		10633 => "11010111",
		10634 => "11111111",
		10635 => "11111111",
		10636 => "11111111",
		10637 => "01001101",
		10638 => "01011001",
		10639 => "11101110",
		10640 => "11111111",
		10641 => "11111111",
		10642 => "11111111",
		10643 => "11111111",
		10644 => "11111111",
		10645 => "11111111",
		10646 => "11111111",
		10647 => "11111111",
		10648 => "11111111",
		10649 => "11111111",
		10650 => "11111111",
		10651 => "11111111",
		10652 => "11011100",
		10653 => "01000111",
		10654 => "10101110",
		10655 => "11111111",
		10656 => "11111111",
		10657 => "11111111",
		10658 => "11111111",
		10659 => "11111111",
		10660 => "01110000",
		10661 => "01000111",
		10662 => "10000001",
		10663 => "11100010",
		10664 => "11101110",
		10665 => "10011000",
		10666 => "01000111",
		10667 => "01110000",
		10668 => "01111100",
		10669 => "10101110",
		10670 => "11111001",
		10671 => "11111111",
		10672 => "11111111",
		10673 => "10101001",
		10674 => "01000111",
		10675 => "01110000",
		10676 => "01010011",
		10677 => "01000111",
		10678 => "11111111",
		10679 => "11111111",
		10680 => "11111111",
		10681 => "11111111",
		10682 => "11111111",
		10683 => "11111111",
		10684 => "11111111",
		10685 => "11111111",
		10686 => "10111010",
		10687 => "01000111",
		10688 => "11011100",
		10689 => "11011100",
		10690 => "01000111",
		10691 => "10111010",
		10692 => "11111111",
		10693 => "11111111",
		10694 => "11111111",
		10695 => "11111111",
		10696 => "11111111",
		10697 => "11111111",
		10698 => "01011001",
		10699 => "01000111",
		10700 => "01110000",
		10701 => "01101010",
		10702 => "01001101",
		10703 => "11110011",
		10704 => "11111111",
		10705 => "11111111",
		10706 => "11101110",
		10707 => "10100011",
		10708 => "01110101",
		10709 => "01011110",
		10710 => "01011001",
		10711 => "11101110",
		10712 => "11111111",
		10713 => "11011100",
		10714 => "01110000",
		10715 => "01000111",
		10716 => "01011001",
		10717 => "11101110",
		10718 => "11111111",
		10719 => "11111111",
		10720 => "11111111",
		10721 => "11111111",
		10722 => "11000101",
		10723 => "01000111",
		10724 => "11000101",
		10725 => "11111111",
		10726 => "11111111",
		10727 => "11111111",
		10728 => "11111111",
		10729 => "11111111",
		10730 => "11111111",
		10731 => "11111111",
		10732 => "11111111",
		10733 => "11111001",
		10734 => "10000111",
		10735 => "11111111",
		10736 => "11111111",
		10737 => "11000101",
		10738 => "10001100",
		10739 => "01000111",
		10740 => "01000111",
		10741 => "01011110",
		10742 => "10011000",
		10743 => "11011100",
		10744 => "11111111",
		10745 => "10101001",
		10746 => "10111010",
		10747 => "11111111",
		10748 => "11111111",
		10749 => "11111111",
		10750 => "11111111",
		10751 => "11111111",
		10752 => "11111111",
		10753 => "11111111",
		10754 => "11111111",
		10755 => "11111111",
		10756 => "11111111",
		10757 => "11111111",
		10758 => "11110011",
		10759 => "01100100",
		10760 => "11111111",
		10761 => "11111111",
		10762 => "11111111",
		10763 => "11111111",
		10764 => "11111111",
		10765 => "01000111",
		10766 => "11000000",
		10767 => "11111111",
		10768 => "11111111",
		10769 => "11111111",
		10770 => "11111111",
		10771 => "11111111",
		10772 => "11111111",
		10773 => "11111111",
		10774 => "11111111",
		10775 => "11111111",
		10776 => "11111111",
		10777 => "11111111",
		10778 => "11111111",
		10779 => "11111111",
		10780 => "11111111",
		10781 => "10000001",
		10782 => "01001101",
		10783 => "11101110",
		10784 => "11111111",
		10785 => "11111111",
		10786 => "11111111",
		10787 => "11111111",
		10788 => "11101000",
		10789 => "01010011",
		10790 => "01000111",
		10791 => "01000111",
		10792 => "01000111",
		10793 => "01000111",
		10794 => "10011000",
		10795 => "11111111",
		10796 => "11111111",
		10797 => "11111111",
		10798 => "11111111",
		10799 => "11111111",
		10800 => "11111111",
		10801 => "11000101",
		10802 => "01000111",
		10803 => "01101010",
		10804 => "10000111",
		10805 => "11000000",
		10806 => "11111111",
		10807 => "11100010",
		10808 => "10101001",
		10809 => "11111001",
		10810 => "11111111",
		10811 => "11111111",
		10812 => "11111111",
		10813 => "11111111",
		10814 => "11000101",
		10815 => "01000111",
		10816 => "11011100",
		10817 => "11101000",
		10818 => "01000111",
		10819 => "10111010",
		10820 => "11111111",
		10821 => "11111111",
		10822 => "11111111",
		10823 => "11110011",
		10824 => "10101110",
		10825 => "11111111",
		10826 => "11101110",
		10827 => "10000111",
		10828 => "01110101",
		10829 => "01011110",
		10830 => "01000111",
		10831 => "11110011",
		10832 => "11111111",
		10833 => "11111111",
		10834 => "11111111",
		10835 => "11111111",
		10836 => "11111111",
		10837 => "11101000",
		10838 => "01011001",
		10839 => "01000111",
		10840 => "01011110",
		10841 => "01000111",
		10842 => "01000111",
		10843 => "01000111",
		10844 => "11000101",
		10845 => "11111111",
		10846 => "11111111",
		10847 => "11111111",
		10848 => "11111111",
		10849 => "11111001",
		10850 => "01011001",
		10851 => "01101010",
		10852 => "11111111",
		10853 => "11111111",
		10854 => "11111111",
		10855 => "11111111",
		10856 => "11111111",
		10857 => "11111111",
		10858 => "11111111",
		10859 => "11111111",
		10860 => "11111111",
		10861 => "11111111",
		10862 => "11111111",
		10863 => "11111111",
		10864 => "11111111",
		10865 => "11111111",
		10866 => "11111111",
		10867 => "11000000",
		10868 => "10000111",
		10869 => "01001101",
		10870 => "01000111",
		10871 => "01000111",
		10872 => "01011110",
		10873 => "01001101",
		10874 => "11111001",
		10875 => "11111111",
		10876 => "11111111",
		10877 => "11111111",
		10878 => "11111111",
		10879 => "11111111",
		10880 => "11111111",
		10881 => "11111111",
		10882 => "11111111",
		10883 => "11111111",
		10884 => "11111111",
		10885 => "11111111",
		10886 => "11111111",
		10887 => "11000000",
		10888 => "11111111",
		10889 => "11111111",
		10890 => "11111111",
		10891 => "11111111",
		10892 => "10110100",
		10893 => "01111100",
		10894 => "11111111",
		10895 => "11111111",
		10896 => "11111111",
		10897 => "11111111",
		10898 => "11111111",
		10899 => "10011000",
		10900 => "11111001",
		10901 => "11111111",
		10902 => "11111111",
		10903 => "11111111",
		10904 => "11111111",
		10905 => "11111111",
		10906 => "11111111",
		10907 => "11111111",
		10908 => "11111111",
		10909 => "11100010",
		10910 => "01001101",
		10911 => "10000111",
		10912 => "11111111",
		10913 => "11111111",
		10914 => "11111111",
		10915 => "11111111",
		10916 => "11111111",
		10917 => "11000101",
		10918 => "01000111",
		10919 => "01100100",
		10920 => "10101110",
		10921 => "11011100",
		10922 => "11111111",
		10923 => "11111111",
		10924 => "11111111",
		10925 => "11111111",
		10926 => "11111111",
		10927 => "11111111",
		10928 => "11111111",
		10929 => "10001100",
		10930 => "01000111",
		10931 => "11110011",
		10932 => "11111111",
		10933 => "11111111",
		10934 => "11111111",
		10935 => "11010111",
		10936 => "01000111",
		10937 => "10001100",
		10938 => "11111111",
		10939 => "11111111",
		10940 => "11111111",
		10941 => "11111001",
		10942 => "01110101",
		10943 => "01011001",
		10944 => "11111001",
		10945 => "11111111",
		10946 => "01101010",
		10947 => "01100100",
		10948 => "11101110",
		10949 => "11111111",
		10950 => "11110011",
		10951 => "01110101",
		10952 => "01011001",
		10953 => "11111111",
		10954 => "11111111",
		10955 => "11111111",
		10956 => "11111111",
		10957 => "11000101",
		10958 => "01000111",
		10959 => "11000000",
		10960 => "11111111",
		10961 => "11111111",
		10962 => "11111111",
		10963 => "11111111",
		10964 => "11111111",
		10965 => "11111111",
		10966 => "11101000",
		10967 => "10111010",
		10968 => "10001100",
		10969 => "01000111",
		10970 => "01000111",
		10971 => "10011000",
		10972 => "11111111",
		10973 => "11111111",
		10974 => "11111111",
		10975 => "11111111",
		10976 => "11111111",
		10977 => "10011110",
		10978 => "01000111",
		10979 => "11010111",
		10980 => "11111111",
		10981 => "11111111",
		10982 => "11111111",
		10983 => "11111111",
		10984 => "11111111",
		10985 => "11111111",
		10986 => "11111111",
		10987 => "11111111",
		10988 => "11111111",
		10989 => "11111111",
		10990 => "11111111",
		10991 => "11111111",
		10992 => "11111111",
		10993 => "11111111",
		10994 => "11111111",
		10995 => "11111111",
		10996 => "11111111",
		10997 => "11111001",
		10998 => "11000000",
		10999 => "10000111",
		11000 => "01001101",
		11001 => "10000111",
		11002 => "11111111",
		11003 => "11111111",
		11004 => "11111111",
		11005 => "11111111",
		11006 => "11111111",
		11007 => "11111111",
		11008 => "11111111",
		11009 => "11111111",
		11010 => "11111111",
		11011 => "11111111",
		11012 => "11111111",
		11013 => "11111111",
		11014 => "11111111",
		11015 => "11111111",
		11016 => "11111111",
		11017 => "11111111",
		11018 => "11111111",
		11019 => "11101110",
		11020 => "01010011",
		11021 => "11101110",
		11022 => "11111111",
		11023 => "11111111",
		11024 => "11111111",
		11025 => "11111111",
		11026 => "11111111",
		11027 => "01110101",
		11028 => "11000101",
		11029 => "11111111",
		11030 => "11111111",
		11031 => "11111111",
		11032 => "11111111",
		11033 => "11111111",
		11034 => "11111111",
		11035 => "11111111",
		11036 => "11111111",
		11037 => "11111111",
		11038 => "10100011",
		11039 => "01000111",
		11040 => "11000000",
		11041 => "11111111",
		11042 => "11111111",
		11043 => "11111111",
		11044 => "11111111",
		11045 => "11111111",
		11046 => "10010011",
		11047 => "01001101",
		11048 => "11010111",
		11049 => "11111111",
		11050 => "11111111",
		11051 => "11111111",
		11052 => "11111111",
		11053 => "11000000",
		11054 => "01100100",
		11055 => "10011000",
		11056 => "01110000",
		11057 => "01000111",
		11058 => "10010011",
		11059 => "11111111",
		11060 => "11111111",
		11061 => "11111111",
		11062 => "11111111",
		11063 => "11111111",
		11064 => "10010011",
		11065 => "01000111",
		11066 => "01011001",
		11067 => "01110101",
		11068 => "01110101",
		11069 => "01011110",
		11070 => "01000111",
		11071 => "11000101",
		11072 => "11111111",
		11073 => "11111111",
		11074 => "11010001",
		11075 => "01010011",
		11076 => "01000111",
		11077 => "01110101",
		11078 => "01000111",
		11079 => "01000111",
		11080 => "11000000",
		11081 => "11111111",
		11082 => "11111111",
		11083 => "11111111",
		11084 => "11111111",
		11085 => "11110011",
		11086 => "01100100",
		11087 => "01010011",
		11088 => "10011110",
		11089 => "10111010",
		11090 => "10110100",
		11091 => "11111111",
		11092 => "11111111",
		11093 => "11111111",
		11094 => "11111111",
		11095 => "11111111",
		11096 => "10101110",
		11097 => "01000111",
		11098 => "01110101",
		11099 => "11111111",
		11100 => "11111111",
		11101 => "11111111",
		11102 => "11111111",
		11103 => "11111111",
		11104 => "11100010",
		11105 => "01001101",
		11106 => "10001100",
		11107 => "11111111",
		11108 => "11111111",
		11109 => "11111111",
		11110 => "11111111",
		11111 => "11111111",
		11112 => "11111111",
		11113 => "11111111",
		11114 => "11111111",
		11115 => "11111111",
		11116 => "11110011",
		11117 => "10001100",
		11118 => "11010001",
		11119 => "11111111",
		11120 => "11111111",
		11121 => "11111111",
		11122 => "11111111",
		11123 => "11111111",
		11124 => "11111111",
		11125 => "11111111",
		11126 => "11111111",
		11127 => "11111111",
		11128 => "10001100",
		11129 => "11000101",
		11130 => "11111111",
		11131 => "11111111",
		11132 => "11111111",
		11133 => "11111111",
		11134 => "11111111",
		11135 => "11111111",
		11136 => "11111111",
		11137 => "11111111",
		11138 => "11111111",
		11139 => "11111111",
		11140 => "11111111",
		11141 => "11111111",
		11142 => "11111111",
		11143 => "11111111",
		11144 => "11111111",
		11145 => "11111111",
		11146 => "11111111",
		11147 => "10000001",
		11148 => "01000111",
		11149 => "11111111",
		11150 => "11111111",
		11151 => "11111111",
		11152 => "11111001",
		11153 => "10111010",
		11154 => "01110101",
		11155 => "01000111",
		11156 => "01111100",
		11157 => "11111111",
		11158 => "11111111",
		11159 => "11111111",
		11160 => "11111111",
		11161 => "11111111",
		11162 => "11111111",
		11163 => "11111111",
		11164 => "11111111",
		11165 => "11111111",
		11166 => "11111001",
		11167 => "01110000",
		11168 => "01011001",
		11169 => "11111111",
		11170 => "11111111",
		11171 => "11111111",
		11172 => "11111111",
		11173 => "11111111",
		11174 => "11111001",
		11175 => "01100100",
		11176 => "01011110",
		11177 => "11110011",
		11178 => "11111111",
		11179 => "11111111",
		11180 => "11111111",
		11181 => "11100010",
		11182 => "01000111",
		11183 => "01000111",
		11184 => "01010011",
		11185 => "10011110",
		11186 => "11111001",
		11187 => "11111111",
		11188 => "11111111",
		11189 => "11111001",
		11190 => "11111001",
		11191 => "11111111",
		11192 => "01111100",
		11193 => "01010011",
		11194 => "01000111",
		11195 => "01000111",
		11196 => "01100100",
		11197 => "10001100",
		11198 => "11010111",
		11199 => "11111111",
		11200 => "11111111",
		11201 => "11111111",
		11202 => "11111111",
		11203 => "11101000",
		11204 => "01111100",
		11205 => "01000111",
		11206 => "01001101",
		11207 => "01000111",
		11208 => "10101110",
		11209 => "11111111",
		11210 => "11010111",
		11211 => "11111111",
		11212 => "11111111",
		11213 => "11111111",
		11214 => "11101000",
		11215 => "01110000",
		11216 => "01000111",
		11217 => "01000111",
		11218 => "01101010",
		11219 => "11111111",
		11220 => "11111111",
		11221 => "11111111",
		11222 => "11111111",
		11223 => "11100010",
		11224 => "01001101",
		11225 => "01011110",
		11226 => "11110011",
		11227 => "11111111",
		11228 => "11111111",
		11229 => "11111111",
		11230 => "11111111",
		11231 => "11111111",
		11232 => "01110000",
		11233 => "01011001",
		11234 => "11101110",
		11235 => "11111111",
		11236 => "11111111",
		11237 => "11111111",
		11238 => "11111111",
		11239 => "11111111",
		11240 => "11111111",
		11241 => "11111111",
		11242 => "11111111",
		11243 => "11111111",
		11244 => "01110101",
		11245 => "01110101",
		11246 => "01001101",
		11247 => "10000111",
		11248 => "11111111",
		11249 => "11111111",
		11250 => "11111111",
		11251 => "11111111",
		11252 => "11111111",
		11253 => "11111111",
		11254 => "11111111",
		11255 => "11111111",
		11256 => "10101110",
		11257 => "11111001",
		11258 => "11111111",
		11259 => "11111111",
		11260 => "11111111",
		11261 => "11111111",
		11262 => "11111111",
		11263 => "11111111",
		11264 => "11111111",
		11265 => "11111111",
		11266 => "11111111",
		11267 => "11111111",
		11268 => "11111111",
		11269 => "11111111",
		11270 => "11111111",
		11271 => "11111111",
		11272 => "11111111",
		11273 => "11111111",
		11274 => "11000101",
		11275 => "01000111",
		11276 => "01110000",
		11277 => "11111111",
		11278 => "11010001",
		11279 => "10001100",
		11280 => "01001101",
		11281 => "01110101",
		11282 => "10111010",
		11283 => "11110011",
		11284 => "01111100",
		11285 => "11101000",
		11286 => "11111111",
		11287 => "11111111",
		11288 => "11111111",
		11289 => "11111111",
		11290 => "11111111",
		11291 => "11111111",
		11292 => "11111111",
		11293 => "11111111",
		11294 => "11111111",
		11295 => "11100010",
		11296 => "01001101",
		11297 => "11111111",
		11298 => "11111111",
		11299 => "11111111",
		11300 => "11111111",
		11301 => "11111111",
		11302 => "11111111",
		11303 => "11011100",
		11304 => "01001101",
		11305 => "10000111",
		11306 => "11111111",
		11307 => "11111111",
		11308 => "11111111",
		11309 => "11111111",
		11310 => "01011001",
		11311 => "01111100",
		11312 => "11111111",
		11313 => "11111111",
		11314 => "11111111",
		11315 => "11111111",
		11316 => "11111111",
		11317 => "11000101",
		11318 => "01011001",
		11319 => "01101010",
		11320 => "01000111",
		11321 => "10101110",
		11322 => "11010111",
		11323 => "01011110",
		11324 => "01010011",
		11325 => "10111010",
		11326 => "11111111",
		11327 => "11111111",
		11328 => "11111111",
		11329 => "11111111",
		11330 => "11111111",
		11331 => "10100011",
		11332 => "01000111",
		11333 => "01101010",
		11334 => "11100010",
		11335 => "01101010",
		11336 => "01000111",
		11337 => "10000001",
		11338 => "01000111",
		11339 => "11110011",
		11340 => "11111111",
		11341 => "11111111",
		11342 => "11111111",
		11343 => "11111111",
		11344 => "11101110",
		11345 => "01000111",
		11346 => "10010011",
		11347 => "11111111",
		11348 => "11111111",
		11349 => "11111111",
		11350 => "11111001",
		11351 => "01100100",
		11352 => "01010011",
		11353 => "11101000",
		11354 => "11111111",
		11355 => "11111111",
		11356 => "11111111",
		11357 => "11111111",
		11358 => "11111111",
		11359 => "10101001",
		11360 => "01000111",
		11361 => "11000000",
		11362 => "11111111",
		11363 => "11111111",
		11364 => "11111111",
		11365 => "11111111",
		11366 => "11111111",
		11367 => "11111111",
		11368 => "11111111",
		11369 => "11111111",
		11370 => "11111111",
		11371 => "10101001",
		11372 => "10010011",
		11373 => "11111111",
		11374 => "11111111",
		11375 => "11111111",
		11376 => "11111111",
		11377 => "11111111",
		11378 => "11111111",
		11379 => "11111111",
		11380 => "11111111",
		11381 => "11111111",
		11382 => "11111111",
		11383 => "11111111",
		11384 => "11111111",
		11385 => "11111111",
		11386 => "11111111",
		11387 => "11111111",
		11388 => "11111111",
		11389 => "11111111",
		11390 => "11111111",
		11391 => "11111111",
		11392 => "11111111",
		11393 => "11111111",
		11394 => "11111111",
		11395 => "11111111",
		11396 => "11111111",
		11397 => "11111111",
		11398 => "11111111",
		11399 => "11111111",
		11400 => "11111111",
		11401 => "11110011",
		11402 => "01011001",
		11403 => "01001101",
		11404 => "11001011",
		11405 => "01011110",
		11406 => "01011110",
		11407 => "10100011",
		11408 => "11101000",
		11409 => "11111111",
		11410 => "11111111",
		11411 => "11111111",
		11412 => "11111111",
		11413 => "11111111",
		11414 => "11111111",
		11415 => "11111111",
		11416 => "11111111",
		11417 => "11111111",
		11418 => "11111111",
		11419 => "11111111",
		11420 => "11111111",
		11421 => "11111111",
		11422 => "11111111",
		11423 => "11111111",
		11424 => "10100011",
		11425 => "11001011",
		11426 => "11111111",
		11427 => "11111111",
		11428 => "11111111",
		11429 => "11111111",
		11430 => "11111111",
		11431 => "11111111",
		11432 => "10101001",
		11433 => "01000111",
		11434 => "10110100",
		11435 => "11111111",
		11436 => "11111111",
		11437 => "11011100",
		11438 => "01000111",
		11439 => "10011000",
		11440 => "11111111",
		11441 => "11111111",
		11442 => "11111111",
		11443 => "11111111",
		11444 => "11111111",
		11445 => "11111001",
		11446 => "01000111",
		11447 => "01000111",
		11448 => "10100011",
		11449 => "11111111",
		11450 => "11111111",
		11451 => "11110011",
		11452 => "10000001",
		11453 => "01000111",
		11454 => "01110000",
		11455 => "11010001",
		11456 => "11111111",
		11457 => "11000101",
		11458 => "01101010",
		11459 => "01000111",
		11460 => "10010011",
		11461 => "11111001",
		11462 => "11111111",
		11463 => "11101110",
		11464 => "01110000",
		11465 => "01000111",
		11466 => "01111100",
		11467 => "11111111",
		11468 => "11111111",
		11469 => "11111111",
		11470 => "11111111",
		11471 => "11111111",
		11472 => "11111111",
		11473 => "01101010",
		11474 => "01011001",
		11475 => "11111111",
		11476 => "11111111",
		11477 => "11111111",
		11478 => "10011000",
		11479 => "01001101",
		11480 => "11010001",
		11481 => "11111111",
		11482 => "11111111",
		11483 => "11111111",
		11484 => "11111111",
		11485 => "11111111",
		11486 => "11101000",
		11487 => "01001101",
		11488 => "10000001",
		11489 => "11111111",
		11490 => "11111111",
		11491 => "11111111",
		11492 => "11111111",
		11493 => "11111111",
		11494 => "11111111",
		11495 => "11111111",
		11496 => "11111111",
		11497 => "11111111",
		11498 => "11111001",
		11499 => "01010011",
		11500 => "11011100",
		11501 => "11111111",
		11502 => "11111111",
		11503 => "11111111",
		11504 => "11111111",
		11505 => "11111111",
		11506 => "11111111",
		11507 => "11111111",
		11508 => "11111111",
		11509 => "11111111",
		11510 => "11111111",
		11511 => "11111111",
		11512 => "11111111",
		11513 => "11111111",
		11514 => "11111111",
		11515 => "11111111",
		11516 => "11111111",
		11517 => "11111111",
		11518 => "11111111",
		11519 => "11111111",
		11520 => "11111111",
		11521 => "11111111",
		11522 => "11111111",
		11523 => "11111111",
		11524 => "11111111",
		11525 => "11111111",
		11526 => "11111111",
		11527 => "11111111",
		11528 => "11111111",
		11529 => "10100011",
		11530 => "01000111",
		11531 => "01001101",
		11532 => "01001101",
		11533 => "11010001",
		11534 => "11111111",
		11535 => "11111111",
		11536 => "11111111",
		11537 => "11111111",
		11538 => "11111111",
		11539 => "11111111",
		11540 => "11111111",
		11541 => "11111111",
		11542 => "10101110",
		11543 => "11111111",
		11544 => "11111111",
		11545 => "11111111",
		11546 => "11111111",
		11547 => "11111111",
		11548 => "11111111",
		11549 => "11111111",
		11550 => "11111111",
		11551 => "11111111",
		11552 => "11111001",
		11553 => "01011001",
		11554 => "11110011",
		11555 => "11111111",
		11556 => "11111111",
		11557 => "11111111",
		11558 => "11111111",
		11559 => "11111111",
		11560 => "11111111",
		11561 => "01111100",
		11562 => "01000111",
		11563 => "01111100",
		11564 => "10010011",
		11565 => "01010011",
		11566 => "01010011",
		11567 => "11101110",
		11568 => "11111111",
		11569 => "11111111",
		11570 => "10111010",
		11571 => "11101110",
		11572 => "11111111",
		11573 => "11101000",
		11574 => "01110101",
		11575 => "01001101",
		11576 => "01011110",
		11577 => "11011100",
		11578 => "11111111",
		11579 => "11111111",
		11580 => "11111111",
		11581 => "11000000",
		11582 => "01011001",
		11583 => "01000111",
		11584 => "01011001",
		11585 => "01000111",
		11586 => "01100100",
		11587 => "11000101",
		11588 => "11111111",
		11589 => "11111111",
		11590 => "11111111",
		11591 => "11000101",
		11592 => "01010011",
		11593 => "01011001",
		11594 => "01101010",
		11595 => "11111111",
		11596 => "11111111",
		11597 => "11111111",
		11598 => "11111111",
		11599 => "11111111",
		11600 => "11111111",
		11601 => "10111010",
		11602 => "01000111",
		11603 => "01110101",
		11604 => "10101110",
		11605 => "01111100",
		11606 => "01000111",
		11607 => "10111010",
		11608 => "11111111",
		11609 => "11111111",
		11610 => "11111111",
		11611 => "11111111",
		11612 => "11111111",
		11613 => "11111111",
		11614 => "01110101",
		11615 => "01010011",
		11616 => "11101110",
		11617 => "11111111",
		11618 => "11111111",
		11619 => "11111111",
		11620 => "11111111",
		11621 => "11111111",
		11622 => "11111111",
		11623 => "11111111",
		11624 => "11111111",
		11625 => "11111111",
		11626 => "11001011",
		11627 => "01010011",
		11628 => "11111111",
		11629 => "11111111",
		11630 => "11111111",
		11631 => "11111111",
		11632 => "11111111",
		11633 => "11010001",
		11634 => "10000111",
		11635 => "01110000",
		11636 => "10101110",
		11637 => "11111111",
		11638 => "11111111",
		11639 => "11111111",
		11640 => "11111111",
		11641 => "11111111",
		11642 => "11111111",
		11643 => "11111111",
		11644 => "11111111",
		11645 => "11111111",
		11646 => "11111111",
		11647 => "11111111",
		11648 => "11111111",
		11649 => "11111111",
		11650 => "11111111",
		11651 => "11111111",
		11652 => "11111111",
		11653 => "11111111",
		11654 => "11111111",
		11655 => "11111111",
		11656 => "11111111",
		11657 => "11010001",
		11658 => "01000111",
		11659 => "10111010",
		11660 => "11111001",
		11661 => "11111111",
		11662 => "11111111",
		11663 => "11111111",
		11664 => "11111111",
		11665 => "11111111",
		11666 => "11111111",
		11667 => "11111111",
		11668 => "11111111",
		11669 => "11111111",
		11670 => "01100100",
		11671 => "11011100",
		11672 => "11111111",
		11673 => "11111111",
		11674 => "11111111",
		11675 => "11111111",
		11676 => "11111111",
		11677 => "11111111",
		11678 => "11111111",
		11679 => "11111111",
		11680 => "11111111",
		11681 => "01001101",
		11682 => "01110101",
		11683 => "11111111",
		11684 => "11111111",
		11685 => "11111111",
		11686 => "11111111",
		11687 => "11111111",
		11688 => "11111111",
		11689 => "11111001",
		11690 => "01110000",
		11691 => "01000111",
		11692 => "01000111",
		11693 => "10000001",
		11694 => "11100010",
		11695 => "11111111",
		11696 => "11111111",
		11697 => "11111001",
		11698 => "01001101",
		11699 => "01011001",
		11700 => "10011000",
		11701 => "01011001",
		11702 => "11101110",
		11703 => "11011100",
		11704 => "01011110",
		11705 => "01001101",
		11706 => "10110100",
		11707 => "11111111",
		11708 => "11110011",
		11709 => "10110100",
		11710 => "01100100",
		11711 => "01000111",
		11712 => "01011110",
		11713 => "10111010",
		11714 => "11111111",
		11715 => "11111111",
		11716 => "11111111",
		11717 => "11111001",
		11718 => "10100011",
		11719 => "01000111",
		11720 => "01101010",
		11721 => "11101110",
		11722 => "01000111",
		11723 => "10000111",
		11724 => "10100011",
		11725 => "10100011",
		11726 => "11111111",
		11727 => "11111111",
		11728 => "11111111",
		11729 => "11111111",
		11730 => "10101110",
		11731 => "01011001",
		11732 => "01000111",
		11733 => "01000111",
		11734 => "10011110",
		11735 => "11111111",
		11736 => "11111111",
		11737 => "11111111",
		11738 => "11111111",
		11739 => "11111111",
		11740 => "11111111",
		11741 => "11111111",
		11742 => "01000111",
		11743 => "10111010",
		11744 => "11111111",
		11745 => "11111111",
		11746 => "11111111",
		11747 => "11111111",
		11748 => "11111111",
		11749 => "11111111",
		11750 => "11111111",
		11751 => "11111111",
		11752 => "11111111",
		11753 => "11111111",
		11754 => "10111010",
		11755 => "01000111",
		11756 => "10111010",
		11757 => "11111111",
		11758 => "11111111",
		11759 => "11011100",
		11760 => "10000001",
		11761 => "01000111",
		11762 => "01000111",
		11763 => "01010011",
		11764 => "01000111",
		11765 => "10101110",
		11766 => "11111111",
		11767 => "11111111",
		11768 => "11111111",
		11769 => "11111111",
		11770 => "11111111",
		11771 => "11111111",
		11772 => "11111111",
		11773 => "11111111",
		11774 => "11111111",
		11775 => "11111111",
		11776 => "11111111",
		11777 => "11111111",
		11778 => "11111111",
		11779 => "11111111",
		11780 => "11111111",
		11781 => "11111111",
		11782 => "11111111",
		11783 => "11111111",
		11784 => "11111111",
		11785 => "11111111",
		11786 => "01011110",
		11787 => "11111111",
		11788 => "11111111",
		11789 => "11111111",
		11790 => "11111111",
		11791 => "11111111",
		11792 => "11111111",
		11793 => "11111111",
		11794 => "11111111",
		11795 => "11111111",
		11796 => "11111111",
		11797 => "11000000",
		11798 => "01010011",
		11799 => "01101010",
		11800 => "11111111",
		11801 => "11111111",
		11802 => "11111111",
		11803 => "11111111",
		11804 => "11111111",
		11805 => "11111111",
		11806 => "11111111",
		11807 => "11111111",
		11808 => "11111111",
		11809 => "10111010",
		11810 => "01000111",
		11811 => "10011000",
		11812 => "11111111",
		11813 => "11111111",
		11814 => "11111111",
		11815 => "11111111",
		11816 => "11111111",
		11817 => "11111111",
		11818 => "11110011",
		11819 => "01100100",
		11820 => "01010011",
		11821 => "11011100",
		11822 => "11111111",
		11823 => "11111111",
		11824 => "11111111",
		11825 => "11111111",
		11826 => "11010111",
		11827 => "01000111",
		11828 => "01000111",
		11829 => "01001101",
		11830 => "11111111",
		11831 => "11111111",
		11832 => "11110011",
		11833 => "01110101",
		11834 => "01000111",
		11835 => "01100100",
		11836 => "01010011",
		11837 => "01000111",
		11838 => "01101010",
		11839 => "10111010",
		11840 => "11111111",
		11841 => "11111111",
		11842 => "11111111",
		11843 => "11111111",
		11844 => "11000101",
		11845 => "01011110",
		11846 => "01000111",
		11847 => "10000001",
		11848 => "11111001",
		11849 => "11111111",
		11850 => "10100011",
		11851 => "01000111",
		11852 => "01000111",
		11853 => "01011001",
		11854 => "11111111",
		11855 => "11111111",
		11856 => "11111111",
		11857 => "11111111",
		11858 => "11111111",
		11859 => "11001011",
		11860 => "01001101",
		11861 => "10000001",
		11862 => "11111111",
		11863 => "11111111",
		11864 => "11111111",
		11865 => "11111111",
		11866 => "11111111",
		11867 => "11111111",
		11868 => "11111111",
		11869 => "11010001",
		11870 => "10000111",
		11871 => "11111111",
		11872 => "11111111",
		11873 => "11111111",
		11874 => "11111111",
		11875 => "11111111",
		11876 => "11111111",
		11877 => "11111111",
		11878 => "11111111",
		11879 => "11111111",
		11880 => "11111111",
		11881 => "11111111",
		11882 => "11101110",
		11883 => "01001101",
		11884 => "01001101",
		11885 => "10000001",
		11886 => "01110101",
		11887 => "01000111",
		11888 => "01000111",
		11889 => "01010011",
		11890 => "10101110",
		11891 => "11111111",
		11892 => "10101110",
		11893 => "01011001",
		11894 => "11111111",
		11895 => "11111111",
		11896 => "11111111",
		11897 => "11111111",
		11898 => "11111111",
		11899 => "11111111",
		11900 => "11111111",
		11901 => "11111111",
		11902 => "11111111",
		11903 => "11111111",
		11904 => "11111111",
		11905 => "11111111",
		11906 => "11111111",
		11907 => "11111111",
		11908 => "11111111",
		11909 => "11111111",
		11910 => "11111111",
		11911 => "11111111",
		11912 => "11111111",
		11913 => "11111111",
		11914 => "11011100",
		11915 => "11111111",
		11916 => "11111111",
		11917 => "11111111",
		11918 => "11111111",
		11919 => "11111111",
		11920 => "11111111",
		11921 => "11111111",
		11922 => "11111111",
		11923 => "11100010",
		11924 => "01111100",
		11925 => "01000111",
		11926 => "01000111",
		11927 => "01011110",
		11928 => "10101001",
		11929 => "11111111",
		11930 => "11111111",
		11931 => "11111111",
		11932 => "11111111",
		11933 => "11111111",
		11934 => "11111111",
		11935 => "11111111",
		11936 => "11111111",
		11937 => "11111111",
		11938 => "10011000",
		11939 => "01000111",
		11940 => "10100011",
		11941 => "11111111",
		11942 => "11111111",
		11943 => "11111111",
		11944 => "11111111",
		11945 => "11111111",
		11946 => "11111111",
		11947 => "11101000",
		11948 => "01011110",
		11949 => "01010011",
		11950 => "11011100",
		11951 => "11111111",
		11952 => "11111111",
		11953 => "11111111",
		11954 => "11111111",
		11955 => "01011110",
		11956 => "01001101",
		11957 => "01000111",
		11958 => "11010111",
		11959 => "11101000",
		11960 => "10101001",
		11961 => "01100100",
		11962 => "01000111",
		11963 => "01001101",
		11964 => "10001100",
		11965 => "11010111",
		11966 => "11111111",
		11967 => "11111111",
		11968 => "11111111",
		11969 => "11111111",
		11970 => "11000101",
		11971 => "01110101",
		11972 => "01000111",
		11973 => "01101010",
		11974 => "11010001",
		11975 => "11111111",
		11976 => "11111111",
		11977 => "11111111",
		11978 => "01100100",
		11979 => "01000111",
		11980 => "01000111",
		11981 => "10011110",
		11982 => "11111111",
		11983 => "11111111",
		11984 => "11111111",
		11985 => "11111111",
		11986 => "11001011",
		11987 => "01001101",
		11988 => "01110000",
		11989 => "11111001",
		11990 => "11111111",
		11991 => "11111111",
		11992 => "11111111",
		11993 => "11111111",
		11994 => "11111111",
		11995 => "11111111",
		11996 => "11011100",
		11997 => "01010011",
		11998 => "11111001",
		11999 => "11111111",
		12000 => "11111111",
		12001 => "11111111",
		12002 => "11111111",
		12003 => "11111111",
		12004 => "11111111",
		12005 => "11111111",
		12006 => "11111111",
		12007 => "11111111",
		12008 => "11111111",
		12009 => "11111111",
		12010 => "11111111",
		12011 => "11000000",
		12012 => "01001101",
		12013 => "01000111",
		12014 => "01000111",
		12015 => "01000111",
		12016 => "10011000",
		12017 => "11110011",
		12018 => "11111111",
		12019 => "11111111",
		12020 => "11110011",
		12021 => "01001101",
		12022 => "11111111",
		12023 => "11111111",
		12024 => "11111111",
		12025 => "11111111",
		12026 => "11111111",
		12027 => "11111111",
		12028 => "11111111",
		12029 => "11111111",
		12030 => "11111111",
		12031 => "11111111",
		12032 => "11111111",
		12033 => "11111111",
		12034 => "11111111",
		12035 => "11111111",
		12036 => "11111111",
		12037 => "11111111",
		12038 => "11111111",
		12039 => "11111111",
		12040 => "11111111",
		12041 => "11111111",
		12042 => "11111111",
		12043 => "11111111",
		12044 => "11111111",
		12045 => "11111111",
		12046 => "11111111",
		12047 => "11111111",
		12048 => "11010111",
		12049 => "01100100",
		12050 => "01000111",
		12051 => "01010011",
		12052 => "10111010",
		12053 => "11111111",
		12054 => "11111111",
		12055 => "11111111",
		12056 => "11111111",
		12057 => "11111111",
		12058 => "11111111",
		12059 => "11111111",
		12060 => "11111111",
		12061 => "11111111",
		12062 => "11111111",
		12063 => "11111111",
		12064 => "11111111",
		12065 => "11111111",
		12066 => "11111111",
		12067 => "11111111",
		12068 => "10001100",
		12069 => "01000111",
		12070 => "10001100",
		12071 => "11110011",
		12072 => "11111111",
		12073 => "11111111",
		12074 => "11111111",
		12075 => "11000000",
		12076 => "01000111",
		12077 => "10010011",
		12078 => "01101010",
		12079 => "01001101",
		12080 => "10001100",
		12081 => "10110100",
		12082 => "01101010",
		12083 => "01000111",
		12084 => "11011100",
		12085 => "11111111",
		12086 => "01011001",
		12087 => "10101001",
		12088 => "11101000",
		12089 => "11111111",
		12090 => "11111111",
		12091 => "11111111",
		12092 => "11111001",
		12093 => "11000000",
		12094 => "10000111",
		12095 => "01001101",
		12096 => "01000111",
		12097 => "01111100",
		12098 => "11000101",
		12099 => "11111111",
		12100 => "11111111",
		12101 => "11111111",
		12102 => "11101110",
		12103 => "10011000",
		12104 => "01001101",
		12105 => "01001101",
		12106 => "11111001",
		12107 => "11111111",
		12108 => "10100011",
		12109 => "01000111",
		12110 => "10010011",
		12111 => "11001011",
		12112 => "10000111",
		12113 => "01000111",
		12114 => "01110101",
		12115 => "01011001",
		12116 => "01111100",
		12117 => "11111111",
		12118 => "11111111",
		12119 => "11111111",
		12120 => "11111111",
		12121 => "11111111",
		12122 => "11011100",
		12123 => "01010011",
		12124 => "01011110",
		12125 => "11101000",
		12126 => "11111111",
		12127 => "11111111",
		12128 => "11111111",
		12129 => "11111111",
		12130 => "11111111",
		12131 => "11111111",
		12132 => "11111111",
		12133 => "11111111",
		12134 => "11111111",
		12135 => "11111111",
		12136 => "11111111",
		12137 => "11111111",
		12138 => "11111111",
		12139 => "11111111",
		12140 => "11111111",
		12141 => "11111111",
		12142 => "11111111",
		12143 => "11111111",
		12144 => "11111111",
		12145 => "11111111",
		12146 => "11111111",
		12147 => "11111111",
		12148 => "01111100",
		12149 => "11010111",
		12150 => "11111111",
		12151 => "11111111",
		12152 => "11111111",
		12153 => "11111111",
		12154 => "11111111",
		12155 => "11111111",
		12156 => "11111111",
		12157 => "11111111",
		12158 => "11111111",
		12159 => "11111111",
		12160 => "11111111",
		12161 => "11111111",
		12162 => "11111111",
		12163 => "11111111",
		12164 => "11111111",
		12165 => "11111111",
		12166 => "11111111",
		12167 => "11111111",
		12168 => "11111111",
		12169 => "11111111",
		12170 => "11111111",
		12171 => "11111111",
		12172 => "11101110",
		12173 => "11111111",
		12174 => "11110011",
		12175 => "10001100",
		12176 => "01000111",
		12177 => "01000111",
		12178 => "10001100",
		12179 => "11110011",
		12180 => "11111111",
		12181 => "11111111",
		12182 => "11111111",
		12183 => "11111111",
		12184 => "11111111",
		12185 => "11111111",
		12186 => "11111111",
		12187 => "11111111",
		12188 => "11111111",
		12189 => "11111111",
		12190 => "11111111",
		12191 => "11111111",
		12192 => "11111111",
		12193 => "11111111",
		12194 => "11111111",
		12195 => "11111111",
		12196 => "11111111",
		12197 => "10100011",
		12198 => "01000111",
		12199 => "01011001",
		12200 => "10010011",
		12201 => "10100011",
		12202 => "10000111",
		12203 => "01001101",
		12204 => "10000001",
		12205 => "11111111",
		12206 => "11111001",
		12207 => "10000111",
		12208 => "01000111",
		12209 => "01000111",
		12210 => "01100100",
		12211 => "11010111",
		12212 => "11111111",
		12213 => "11101000",
		12214 => "10100011",
		12215 => "11111111",
		12216 => "11100010",
		12217 => "11000000",
		12218 => "10011110",
		12219 => "01110101",
		12220 => "01001101",
		12221 => "01000111",
		12222 => "01011110",
		12223 => "10011000",
		12224 => "11101000",
		12225 => "11111111",
		12226 => "11111111",
		12227 => "11111111",
		12228 => "11110011",
		12229 => "10011110",
		12230 => "01001101",
		12231 => "01001101",
		12232 => "10011000",
		12233 => "11101110",
		12234 => "11111111",
		12235 => "11111111",
		12236 => "11111001",
		12237 => "10100011",
		12238 => "01001101",
		12239 => "01000111",
		12240 => "01000111",
		12241 => "10010011",
		12242 => "11111111",
		12243 => "10011110",
		12244 => "01000111",
		12245 => "10011110",
		12246 => "11111001",
		12247 => "11111111",
		12248 => "11110011",
		12249 => "10101001",
		12250 => "01010011",
		12251 => "01011110",
		12252 => "11101000",
		12253 => "11111111",
		12254 => "11111111",
		12255 => "11111111",
		12256 => "11111111",
		12257 => "11111111",
		12258 => "11111111",
		12259 => "11111111",
		12260 => "11111111",
		12261 => "11111111",
		12262 => "11111111",
		12263 => "11111111",
		12264 => "11111111",
		12265 => "11111111",
		12266 => "11111111",
		12267 => "11111111",
		12268 => "11111111",
		12269 => "11111111",
		12270 => "11111111",
		12271 => "11111111",
		12272 => "11111111",
		12273 => "11111111",
		12274 => "01111100",
		12275 => "01110000",
		12276 => "10011110",
		12277 => "11111111",
		12278 => "11111111",
		12279 => "11111111",
		12280 => "11111111",
		12281 => "11111111",
		12282 => "11111111",
		12283 => "11111111",
		12284 => "11111111",
		12285 => "11111111",
		12286 => "11111111",
		12287 => "11111111",
		12288 => "11111111",
		12289 => "11111111",
		12290 => "11111111",
		12291 => "11111111",
		12292 => "11111111",
		12293 => "11111111",
		12294 => "11111111",
		12295 => "11111111",
		12296 => "11111111",
		12297 => "11111111",
		12298 => "11111111",
		12299 => "11111111",
		12300 => "11110011",
		12301 => "10011000",
		12302 => "01010011",
		12303 => "01000111",
		12304 => "01100100",
		12305 => "11010111",
		12306 => "11111111",
		12307 => "11111111",
		12308 => "11111111",
		12309 => "11111111",
		12310 => "11111111",
		12311 => "11111111",
		12312 => "11111111",
		12313 => "11111111",
		12314 => "11111111",
		12315 => "11111111",
		12316 => "11111111",
		12317 => "11111111",
		12318 => "11111111",
		12319 => "11111111",
		12320 => "11111111",
		12321 => "11111111",
		12322 => "11111111",
		12323 => "11111111",
		12324 => "11111111",
		12325 => "11111111",
		12326 => "11010111",
		12327 => "10001100",
		12328 => "01001101",
		12329 => "01000111",
		12330 => "01011110",
		12331 => "10101001",
		12332 => "11111001",
		12333 => "11111111",
		12334 => "11111111",
		12335 => "11111111",
		12336 => "10101001",
		12337 => "01000111",
		12338 => "01110000",
		12339 => "11100010",
		12340 => "11000101",
		12341 => "10100011",
		12342 => "01001101",
		12343 => "01001101",
		12344 => "01000111",
		12345 => "01000111",
		12346 => "01000111",
		12347 => "01110101",
		12348 => "10101110",
		12349 => "11100010",
		12350 => "11111111",
		12351 => "11111111",
		12352 => "11111111",
		12353 => "11111111",
		12354 => "11100010",
		12355 => "10011110",
		12356 => "01010011",
		12357 => "01000111",
		12358 => "10001100",
		12359 => "11101110",
		12360 => "11111111",
		12361 => "11111111",
		12362 => "11111111",
		12363 => "11111111",
		12364 => "11111111",
		12365 => "11010111",
		12366 => "01100100",
		12367 => "01001101",
		12368 => "10110100",
		12369 => "11111111",
		12370 => "11111111",
		12371 => "11111111",
		12372 => "10000001",
		12373 => "01000111",
		12374 => "01000111",
		12375 => "01110000",
		12376 => "01001101",
		12377 => "01000111",
		12378 => "10000001",
		12379 => "11110011",
		12380 => "11111111",
		12381 => "11111111",
		12382 => "11111111",
		12383 => "11111111",
		12384 => "11111111",
		12385 => "11111111",
		12386 => "11111111",
		12387 => "11111111",
		12388 => "11111111",
		12389 => "11111111",
		12390 => "11111111",
		12391 => "11111111",
		12392 => "11111111",
		12393 => "11111111",
		12394 => "11111111",
		12395 => "11111111",
		12396 => "11111111",
		12397 => "11111111",
		12398 => "11111111",
		12399 => "11111111",
		12400 => "11111111",
		12401 => "11111111",
		12402 => "11111111",
		12403 => "10011110",
		12404 => "11111111",
		12405 => "11111111",
		12406 => "11111111",
		12407 => "11111111",
		12408 => "11111111",
		12409 => "11111111",
		12410 => "11111111",
		12411 => "11111111",
		12412 => "11111111",
		12413 => "11111111",
		12414 => "11111111",
		12415 => "11111111",
		12416 => "11111111",
		12417 => "11111111",
		12418 => "11111111",
		12419 => "11111111",
		12420 => "11111111",
		12421 => "11111111",
		12422 => "11111111",
		12423 => "11111111",
		12424 => "11111111",
		12425 => "11111111",
		12426 => "11111111",
		12427 => "11111111",
		12428 => "11111111",
		12429 => "01000111",
		12430 => "01001101",
		12431 => "10101001",
		12432 => "11111111",
		12433 => "11111111",
		12434 => "11111111",
		12435 => "11111111",
		12436 => "11111111",
		12437 => "11111111",
		12438 => "11111111",
		12439 => "11111111",
		12440 => "11111111",
		12441 => "11111111",
		12442 => "11111111",
		12443 => "11111111",
		12444 => "11111111",
		12445 => "11111111",
		12446 => "11111111",
		12447 => "11111111",
		12448 => "11111111",
		12449 => "11111111",
		12450 => "11111111",
		12451 => "11111111",
		12452 => "11111111",
		12453 => "11111111",
		12454 => "11111111",
		12455 => "11111111",
		12456 => "11111111",
		12457 => "11111111",
		12458 => "11111111",
		12459 => "11111111",
		12460 => "11111111",
		12461 => "11111111",
		12462 => "11111111",
		12463 => "11111111",
		12464 => "11111111",
		12465 => "11000101",
		12466 => "01010011",
		12467 => "01000111",
		12468 => "01000111",
		12469 => "01000111",
		12470 => "01111100",
		12471 => "10100011",
		12472 => "10111010",
		12473 => "11010001",
		12474 => "11110011",
		12475 => "11111111",
		12476 => "11111111",
		12477 => "11111111",
		12478 => "11111111",
		12479 => "11110011",
		12480 => "10110100",
		12481 => "01101010",
		12482 => "01000111",
		12483 => "01000111",
		12484 => "10001100",
		12485 => "11101000",
		12486 => "11111111",
		12487 => "11111111",
		12488 => "11111111",
		12489 => "11111111",
		12490 => "11111111",
		12491 => "11111001",
		12492 => "10011110",
		12493 => "01000111",
		12494 => "01011001",
		12495 => "11010111",
		12496 => "11111111",
		12497 => "11111111",
		12498 => "11111111",
		12499 => "11111111",
		12500 => "11111111",
		12501 => "11010111",
		12502 => "10100011",
		12503 => "10100011",
		12504 => "10100011",
		12505 => "11011100",
		12506 => "11111111",
		12507 => "11111111",
		12508 => "11111111",
		12509 => "11111111",
		12510 => "11111111",
		12511 => "11111111",
		12512 => "11111111",
		12513 => "11111111",
		12514 => "11111111",
		12515 => "11111111",
		12516 => "11111111",
		12517 => "11111111",
		12518 => "11111111",
		12519 => "11111111",
		12520 => "11111111",
		12521 => "11111111",
		12522 => "11111111",
		12523 => "11111111",
		12524 => "11111111",
		12525 => "11111111",
		12526 => "11111111",
		12527 => "11111111",
		12528 => "11111111",
		12529 => "11111111",
		12530 => "11111111",
		12531 => "11111111",
		12532 => "11111111",
		12533 => "11111111",
		12534 => "11111111",
		12535 => "11111111",
		12536 => "11111111",
		12537 => "11111111",
		12538 => "11111111",
		12539 => "11111111",
		12540 => "11111111",
		12541 => "11111111",
		12542 => "11111111",
		12543 => "11111111",
		12544 => "11111111",
		12545 => "11111111",
		12546 => "11111111",
		12547 => "11111111",
		12548 => "11111111",
		12549 => "11111111",
		12550 => "11111111",
		12551 => "11111111",
		12552 => "11111111",
		12553 => "11111111",
		12554 => "11111111",
		12555 => "11111111",
		12556 => "11111111",
		12557 => "10000111",
		12558 => "10100011",
		12559 => "11111111",
		12560 => "11111111",
		12561 => "11111111",
		12562 => "11111111",
		12563 => "11111111",
		12564 => "11111111",
		12565 => "11111111",
		12566 => "11111111",
		12567 => "11111111",
		12568 => "11111111",
		12569 => "11111111",
		12570 => "11111111",
		12571 => "11111111",
		12572 => "11111111",
		12573 => "11111111",
		12574 => "11111111",
		12575 => "11111111",
		12576 => "11111111",
		12577 => "11111111",
		12578 => "11111111",
		12579 => "11111111",
		12580 => "11111111",
		12581 => "11111111",
		12582 => "11111111",
		12583 => "11111111",
		12584 => "11111111",
		12585 => "11111111",
		12586 => "11111111",
		12587 => "11111111",
		12588 => "11111111",
		12589 => "11111111",
		12590 => "11111111",
		12591 => "11111111",
		12592 => "11111111",
		12593 => "11111111",
		12594 => "01110000",
		12595 => "01011001",
		12596 => "11100010",
		12597 => "11111111",
		12598 => "11111111",
		12599 => "11111111",
		12600 => "11111111",
		12601 => "11111111",
		12602 => "11111111",
		12603 => "11111111",
		12604 => "11101000",
		12605 => "10111010",
		12606 => "10000111",
		12607 => "01000111",
		12608 => "01000111",
		12609 => "01110101",
		12610 => "10111010",
		12611 => "11110011",
		12612 => "11111111",
		12613 => "11111111",
		12614 => "11111111",
		12615 => "11111111",
		12616 => "11111111",
		12617 => "11111111",
		12618 => "11100010",
		12619 => "01101010",
		12620 => "01000111",
		12621 => "01000111",
		12622 => "10011000",
		12623 => "11111111",
		12624 => "11111111",
		12625 => "11111111",
		12626 => "11111111",
		12627 => "11111111",
		12628 => "11111111",
		12629 => "11111111",
		12630 => "11111111",
		12631 => "11111111",
		12632 => "11111111",
		12633 => "11111111",
		12634 => "11111111",
		12635 => "11111111",
		12636 => "11111111",
		12637 => "11111111",
		12638 => "11111111",
		12639 => "11111111",
		12640 => "11111111",
		12641 => "11111111",
		12642 => "11111111",
		12643 => "11111111",
		12644 => "11111111",
		12645 => "11111111",
		12646 => "11111111",
		12647 => "11111111",
		12648 => "11111111",
		12649 => "11111111",
		12650 => "11111111",
		12651 => "11111111",
		12652 => "11111111",
		12653 => "11111111",
		12654 => "11111111",
		12655 => "11111111",
		12656 => "11111111",
		12657 => "11111111",
		12658 => "11111111",
		12659 => "11111111",
		12660 => "11111111",
		12661 => "11111111",
		12662 => "11111111",
		12663 => "11111111",
		12664 => "11111111",
		12665 => "11111111",
		12666 => "11111111",
		12667 => "11111111",
		12668 => "11111111",
		12669 => "11111111",
		12670 => "11111111",
		12671 => "11111111",
		12672 => "11111111",
		12673 => "11111111",
		12674 => "11111111",
		12675 => "11111111",
		12676 => "11111111",
		12677 => "11111111",
		12678 => "11111111",
		12679 => "11111111",
		12680 => "11111111",
		12681 => "11111111",
		12682 => "11111111",
		12683 => "11111111",
		12684 => "11111111",
		12685 => "11101110",
		12686 => "10011110",
		12687 => "11111111",
		12688 => "11111111",
		12689 => "11111111",
		12690 => "11111111",
		12691 => "11111111",
		12692 => "11111111",
		12693 => "11111111",
		12694 => "11111111",
		12695 => "11111111",
		12696 => "11111111",
		12697 => "11111111",
		12698 => "11111111",
		12699 => "11111111",
		12700 => "11111111",
		12701 => "11111111",
		12702 => "11111111",
		12703 => "11111111",
		12704 => "11111111",
		12705 => "11111111",
		12706 => "11111111",
		12707 => "11111111",
		12708 => "11111111",
		12709 => "11111111",
		12710 => "11111111",
		12711 => "11111111",
		12712 => "11111111",
		12713 => "11111111",
		12714 => "11111111",
		12715 => "11111111",
		12716 => "11111111",
		12717 => "11111111",
		12718 => "11111111",
		12719 => "11111111",
		12720 => "11111111",
		12721 => "11111111",
		12722 => "01000111",
		12723 => "10011000",
		12724 => "11111111",
		12725 => "11111111",
		12726 => "11111111",
		12727 => "11111111",
		12728 => "11010111",
		12729 => "10101110",
		12730 => "10000001",
		12731 => "01011001",
		12732 => "01000111",
		12733 => "01000111",
		12734 => "01101010",
		12735 => "10101110",
		12736 => "11101110",
		12737 => "11111111",
		12738 => "11111111",
		12739 => "11111111",
		12740 => "11111111",
		12741 => "11111111",
		12742 => "11111111",
		12743 => "11111111",
		12744 => "11111111",
		12745 => "11110011",
		12746 => "01001101",
		12747 => "01010011",
		12748 => "10111010",
		12749 => "01100100",
		12750 => "01111100",
		12751 => "11111111",
		12752 => "11111111",
		12753 => "11111111",
		12754 => "11111111",
		12755 => "11111111",
		12756 => "11111111",
		12757 => "11111111",
		12758 => "11111111",
		12759 => "11111111",
		12760 => "11111111",
		12761 => "11111111",
		12762 => "11111111",
		12763 => "11111111",
		12764 => "11111111",
		12765 => "11111111",
		12766 => "11111111",
		12767 => "11111111",
		12768 => "11111111",
		12769 => "11111111",
		12770 => "11111111",
		12771 => "11111111",
		12772 => "11111111",
		12773 => "11111111",
		12774 => "11111111",
		12775 => "11111111",
		12776 => "11111111",
		12777 => "11111111",
		12778 => "11111111",
		12779 => "11111111",
		12780 => "11111111",
		12781 => "11111111",
		12782 => "11111111",
		12783 => "11111111",
		12784 => "11111111",
		12785 => "11111111",
		12786 => "11111111",
		12787 => "11111111",
		12788 => "11111111",
		12789 => "11111111",
		12790 => "11111111",
		12791 => "11111111",
		12792 => "11111111",
		12793 => "11111111",
		12794 => "11111111",
		12795 => "11111111",
		12796 => "11111111",
		12797 => "11111111",
		12798 => "11111111",
		12799 => "11111111",
		12800 => "11111111",
		12801 => "11111111",
		12802 => "11111111",
		12803 => "11111111",
		12804 => "11111111",
		12805 => "11111111",
		12806 => "11111111",
		12807 => "11111111",
		12808 => "11111111",
		12809 => "11111111",
		12810 => "11111111",
		12811 => "11111111",
		12812 => "11111111",
		12813 => "11111111",
		12814 => "11111111",
		12815 => "11111111",
		12816 => "11111111",
		12817 => "11111111",
		12818 => "11111111",
		12819 => "11111111",
		12820 => "11111111",
		12821 => "11111111",
		12822 => "11111111",
		12823 => "11111111",
		12824 => "11111111",
		12825 => "11111111",
		12826 => "11111111",
		12827 => "11111111",
		12828 => "11111111",
		12829 => "11111111",
		12830 => "11111111",
		12831 => "11111111",
		12832 => "11111111",
		12833 => "11111111",
		12834 => "11111111",
		12835 => "11111111",
		12836 => "11111111",
		12837 => "11111111",
		12838 => "11111111",
		12839 => "11111111",
		12840 => "11111111",
		12841 => "11111111",
		12842 => "11111111",
		12843 => "11111111",
		12844 => "11111111",
		12845 => "11111111",
		12846 => "11111111",
		12847 => "11111001",
		12848 => "10110100",
		12849 => "10100011",
		12850 => "01010011",
		12851 => "01011001",
		12852 => "10100011",
		12853 => "01110101",
		12854 => "01001101",
		12855 => "01000111",
		12856 => "01000111",
		12857 => "01000111",
		12858 => "01101010",
		12859 => "10010011",
		12860 => "11000000",
		12861 => "11101110",
		12862 => "11111111",
		12863 => "11111111",
		12864 => "11111111",
		12865 => "11111111",
		12866 => "11111111",
		12867 => "11111111",
		12868 => "11111111",
		12869 => "11111111",
		12870 => "11111111",
		12871 => "11111111",
		12872 => "10101110",
		12873 => "01011001",
		12874 => "01000111",
		12875 => "01100100",
		12876 => "01110000",
		12877 => "01000111",
		12878 => "01101010",
		12879 => "10100011",
		12880 => "10101110",
		12881 => "11111001",
		12882 => "11111111",
		12883 => "11111111",
		12884 => "11111111",
		12885 => "11111111",
		12886 => "11111111",
		12887 => "11111111",
		12888 => "11111111",
		12889 => "11111111",
		12890 => "11111111",
		12891 => "11111111",
		12892 => "11111111",
		12893 => "11111111",
		12894 => "11111111",
		12895 => "11111111",
		12896 => "11111111",
		12897 => "11111111",
		12898 => "11111111",
		12899 => "11111111",
		12900 => "11111111",
		12901 => "11111111",
		12902 => "11111111",
		12903 => "11111111",
		12904 => "11111111",
		12905 => "11111111",
		12906 => "11111111",
		12907 => "11111111",
		12908 => "11111111",
		12909 => "11111111",
		12910 => "11111111",
		12911 => "11111111",
		12912 => "11111111",
		12913 => "11111111",
		12914 => "11111111",
		12915 => "11111111",
		12916 => "11111111",
		12917 => "11111111",
		12918 => "11111111",
		12919 => "11111111",
		12920 => "11111111",
		12921 => "11111111",
		12922 => "11111111",
		12923 => "11111111",
		12924 => "11111111",
		12925 => "11111111",
		12926 => "11111111",
		12927 => "11111111",
		12928 => "11111111",
		12929 => "11111111",
		12930 => "11111111",
		12931 => "11111111",
		12932 => "11111111",
		12933 => "11111111",
		12934 => "11111111",
		12935 => "11111111",
		12936 => "11111111",
		12937 => "11111111",
		12938 => "11111111",
		12939 => "11111111",
		12940 => "11111111",
		12941 => "11111111",
		12942 => "11111111",
		12943 => "11111111",
		12944 => "11111111",
		12945 => "11111111",
		12946 => "11111111",
		12947 => "11111111",
		12948 => "11111111",
		12949 => "11111111",
		12950 => "11111111",
		12951 => "11111111",
		12952 => "11111111",
		12953 => "11111111",
		12954 => "11111111",
		12955 => "11111111",
		12956 => "11111111",
		12957 => "11111111",
		12958 => "11111111",
		12959 => "11111111",
		12960 => "11111111",
		12961 => "11111111",
		12962 => "11111111",
		12963 => "11111111",
		12964 => "11111111",
		12965 => "11111111",
		12966 => "11111111",
		12967 => "11111111",
		12968 => "11111111",
		12969 => "11111111",
		12970 => "11111111",
		12971 => "11111111",
		12972 => "11111111",
		12973 => "11111111",
		12974 => "11001011",
		12975 => "01011110",
		12976 => "01000111",
		12977 => "01000111",
		12978 => "01000111",
		12979 => "01000111",
		12980 => "01010011",
		12981 => "01110101",
		12982 => "10011110",
		12983 => "10100011",
		12984 => "11000101",
		12985 => "11110011",
		12986 => "11111111",
		12987 => "11111111",
		12988 => "11111111",
		12989 => "11111111",
		12990 => "11111111",
		12991 => "11111111",
		12992 => "11111111",
		12993 => "11111111",
		12994 => "11111111",
		12995 => "11111111",
		12996 => "11111111",
		12997 => "11111111",
		12998 => "11000101",
		12999 => "01100100",
		13000 => "01000111",
		13001 => "01110101",
		13002 => "10000111",
		13003 => "01110101",
		13004 => "01110101",
		13005 => "01000111",
		13006 => "01000111",
		13007 => "01000111",
		13008 => "01000111",
		13009 => "01100100",
		13010 => "11010001",
		13011 => "11111111",
		13012 => "11111111",
		13013 => "11111111",
		13014 => "11111111",
		13015 => "11111111",
		13016 => "11111111",
		13017 => "11111111",
		13018 => "11111111",
		13019 => "11111111",
		13020 => "11111111",
		13021 => "11111111",
		13022 => "11111111",
		13023 => "11111111",
		13024 => "11111111",
		13025 => "11111111",
		13026 => "11111111",
		13027 => "11111111",
		13028 => "11111111",
		13029 => "11111111",
		13030 => "11111111",
		13031 => "11111111",
		13032 => "11111111",
		13033 => "11111111",
		13034 => "11111111",
		13035 => "11111111",
		13036 => "11111111",
		13037 => "11111111",
		13038 => "11111111",
		13039 => "11111111",
		13040 => "11111111",
		13041 => "11111111",
		13042 => "11111111",
		13043 => "11111111",
		13044 => "11111111",
		13045 => "11111111",
		13046 => "11111111",
		13047 => "11111111",
		13048 => "11111111",
		13049 => "11111111",
		13050 => "11111111",
		13051 => "11111111",
		13052 => "11111111",
		13053 => "11111111",
		13054 => "11111111",
		13055 => "11111111",
		13056 => "11111111",
		13057 => "11111111",
		13058 => "11111111",
		13059 => "11111111",
		13060 => "11111111",
		13061 => "11111111",
		13062 => "11111111",
		13063 => "11111111",
		13064 => "11111111",
		13065 => "11111111",
		13066 => "11111111",
		13067 => "11111111",
		13068 => "11111111",
		13069 => "11111111",
		13070 => "11111111",
		13071 => "11111111",
		13072 => "11111111",
		13073 => "11111111",
		13074 => "11111111",
		13075 => "11111111",
		13076 => "11111111",
		13077 => "11111111",
		13078 => "11111111",
		13079 => "11111111",
		13080 => "11111111",
		13081 => "11111111",
		13082 => "11111111",
		13083 => "11111111",
		13084 => "11111111",
		13085 => "11111111",
		13086 => "11111111",
		13087 => "11111111",
		13088 => "11111111",
		13089 => "11111111",
		13090 => "11111111",
		13091 => "11111111",
		13092 => "11111111",
		13093 => "11111111",
		13094 => "11111111",
		13095 => "11111111",
		13096 => "11111111",
		13097 => "11111111",
		13098 => "11111111",
		13099 => "11111111",
		13100 => "11111111",
		13101 => "11011100",
		13102 => "01001101",
		13103 => "01110101",
		13104 => "11011100",
		13105 => "11111111",
		13106 => "11111111",
		13107 => "11111111",
		13108 => "11111111",
		13109 => "11111111",
		13110 => "11111111",
		13111 => "11111111",
		13112 => "11111111",
		13113 => "11111111",
		13114 => "11111111",
		13115 => "11111111",
		13116 => "11111111",
		13117 => "11111111",
		13118 => "11111111",
		13119 => "11111111",
		13120 => "11111111",
		13121 => "11111111",
		13122 => "11111111",
		13123 => "11111111",
		13124 => "11000000",
		13125 => "01110101",
		13126 => "01000111",
		13127 => "01110101",
		13128 => "11010001",
		13129 => "11111111",
		13130 => "11111111",
		13131 => "11111111",
		13132 => "11111111",
		13133 => "11111111",
		13134 => "11111111",
		13135 => "11111111",
		13136 => "11011100",
		13137 => "01101010",
		13138 => "01011001",
		13139 => "11111001",
		13140 => "11111111",
		13141 => "11111111",
		13142 => "11111111",
		13143 => "11111111",
		13144 => "11111111",
		13145 => "11111111",
		13146 => "11111111",
		13147 => "11111111",
		13148 => "11111111",
		13149 => "11111111",
		13150 => "11111111",
		13151 => "11111111",
		13152 => "11111111",
		13153 => "11111111",
		13154 => "11111111",
		13155 => "11111111",
		13156 => "11111111",
		13157 => "11111111",
		13158 => "11111111",
		13159 => "11111111",
		13160 => "11111111",
		13161 => "11111111",
		13162 => "11111111",
		13163 => "11111111",
		13164 => "11111111",
		13165 => "11111111",
		13166 => "11111111",
		13167 => "11111111",
		13168 => "11111111",
		13169 => "11111111",
		13170 => "11111111",
		13171 => "11111111",
		13172 => "11111111",
		13173 => "11111111",
		13174 => "11111111",
		13175 => "11111111",
		13176 => "11111111",
		13177 => "11111111",
		13178 => "11111111",
		13179 => "11111111",
		13180 => "11111111",
		13181 => "11111111",
		13182 => "11111111",
		13183 => "11111111",
		13184 => "11111111",
		13185 => "11111111",
		13186 => "11111111",
		13187 => "11111111",
		13188 => "11111111",
		13189 => "11111111",
		13190 => "11111111",
		13191 => "11111111",
		13192 => "11111111",
		13193 => "11111111",
		13194 => "11111111",
		13195 => "11111111",
		13196 => "11111111",
		13197 => "11111111",
		13198 => "11111111",
		13199 => "11111111",
		13200 => "11111111",
		13201 => "11111111",
		13202 => "11111111",
		13203 => "11111111",
		13204 => "11111111",
		13205 => "11111111",
		13206 => "11111111",
		13207 => "11111111",
		13208 => "11111111",
		13209 => "11111111",
		13210 => "11111111",
		13211 => "11111111",
		13212 => "11111111",
		13213 => "11111111",
		13214 => "11111111",
		13215 => "11111111",
		13216 => "11111111",
		13217 => "11111111",
		13218 => "11111111",
		13219 => "11111111",
		13220 => "11111111",
		13221 => "11111111",
		13222 => "11111111",
		13223 => "11111111",
		13224 => "11111111",
		13225 => "11111111",
		13226 => "11111111",
		13227 => "11111111",
		13228 => "11111111",
		13229 => "10101001",
		13230 => "01000111",
		13231 => "11110011",
		13232 => "11111111",
		13233 => "11111111",
		13234 => "11111111",
		13235 => "11111111",
		13236 => "11111111",
		13237 => "11111111",
		13238 => "11111111",
		13239 => "11111111",
		13240 => "11111111",
		13241 => "11111111",
		13242 => "11111111",
		13243 => "11111111",
		13244 => "11111111",
		13245 => "11111111",
		13246 => "11111111",
		13247 => "11111111",
		13248 => "11111111",
		13249 => "11101000",
		13250 => "10011110",
		13251 => "01011001",
		13252 => "01000111",
		13253 => "01110101",
		13254 => "11010001",
		13255 => "11111111",
		13256 => "11111111",
		13257 => "11111111",
		13258 => "11111111",
		13259 => "11111111",
		13260 => "11111111",
		13261 => "11111111",
		13262 => "11111111",
		13263 => "11111111",
		13264 => "11111111",
		13265 => "11001011",
		13266 => "01000111",
		13267 => "11010001",
		13268 => "11111111",
		13269 => "11111111",
		13270 => "11111111",
		13271 => "11111111",
		13272 => "11111111",
		13273 => "11111111",
		13274 => "11111111",
		13275 => "11111111",
		13276 => "11111111",
		13277 => "11111111",
		13278 => "11111111",
		13279 => "11111111",
		13280 => "11111111",
		13281 => "11111111",
		13282 => "11111111",
		13283 => "11111111",
		13284 => "11110011",
		13285 => "11101110",
		13286 => "11111111",
		13287 => "11111111",
		13288 => "11111111",
		13289 => "11111111",
		13290 => "11111111",
		13291 => "11111111",
		13292 => "11111111",
		13293 => "11111111",
		13294 => "11111111",
		13295 => "11111111",
		13296 => "11111111",
		13297 => "11111111",
		13298 => "11111111",
		13299 => "11111111",
		13300 => "11111111",
		13301 => "11111111",
		13302 => "11111111",
		13303 => "11111111",
		13304 => "11111111",
		13305 => "11111111",
		13306 => "11111111",
		13307 => "11111111",
		13308 => "11111111",
		13309 => "11111111",
		13310 => "11111111",
		13311 => "11111111",
		13312 => "11111111",
		13313 => "11111111",
		13314 => "11111111",
		13315 => "11111111",
		13316 => "11111111",
		13317 => "11111111",
		13318 => "11111111",
		13319 => "11111111",
		13320 => "11111111",
		13321 => "11111111",
		13322 => "11111111",
		13323 => "11111111",
		13324 => "11111111",
		13325 => "11111111",
		13326 => "11111111",
		13327 => "11111111",
		13328 => "11111111",
		13329 => "11111111",
		13330 => "11111111",
		13331 => "11111111",
		13332 => "11111111",
		13333 => "11111111",
		13334 => "11111111",
		13335 => "11111111",
		13336 => "11111111",
		13337 => "11111111",
		13338 => "11111111",
		13339 => "11111111",
		13340 => "11111111",
		13341 => "11111111",
		13342 => "11111111",
		13343 => "11111111",
		13344 => "11111111",
		13345 => "11111111",
		13346 => "11111111",
		13347 => "11111111",
		13348 => "11111111",
		13349 => "11111111",
		13350 => "11111111",
		13351 => "11111111",
		13352 => "11111111",
		13353 => "11111111",
		13354 => "11111111",
		13355 => "11111111",
		13356 => "11111111",
		13357 => "10101110",
		13358 => "01000111",
		13359 => "11100010",
		13360 => "11111111",
		13361 => "11111111",
		13362 => "11111111",
		13363 => "11111111",
		13364 => "11111111",
		13365 => "11111111",
		13366 => "11111111",
		13367 => "11111111",
		13368 => "11111111",
		13369 => "11111111",
		13370 => "11111111",
		13371 => "11111111",
		13372 => "11111111",
		13373 => "11111111",
		13374 => "11101000",
		13375 => "10110100",
		13376 => "01111100",
		13377 => "01000111",
		13378 => "01000111",
		13379 => "01111100",
		13380 => "11010001",
		13381 => "11111111",
		13382 => "11111111",
		13383 => "11111111",
		13384 => "11111111",
		13385 => "11111111",
		13386 => "11111111",
		13387 => "11111111",
		13388 => "11111111",
		13389 => "11111111",
		13390 => "11111111",
		13391 => "11111111",
		13392 => "11111111",
		13393 => "10101001",
		13394 => "01000111",
		13395 => "11101000",
		13396 => "11111111",
		13397 => "11111111",
		13398 => "11111111",
		13399 => "11111111",
		13400 => "11111111",
		13401 => "11111111",
		13402 => "11111111",
		13403 => "11111111",
		13404 => "11111111",
		13405 => "11111111",
		13406 => "11111111",
		13407 => "11111111",
		13408 => "11111111",
		13409 => "11111111",
		13410 => "11111001",
		13411 => "10000001",
		13412 => "01000111",
		13413 => "01000111",
		13414 => "10001100",
		13415 => "11111001",
		13416 => "11111111",
		13417 => "11111111",
		13418 => "11111111",
		13419 => "11111111",
		13420 => "11111111",
		13421 => "11111111",
		13422 => "11111111",
		13423 => "11111111",
		13424 => "11111111",
		13425 => "11111111",
		13426 => "11111111",
		13427 => "11111111",
		13428 => "11111111",
		13429 => "11111111",
		13430 => "11111111",
		13431 => "11111111",
		13432 => "11111111",
		13433 => "11111111",
		13434 => "11111111",
		13435 => "11111111",
		13436 => "11111111",
		13437 => "11111111",
		13438 => "11111111",
		13439 => "11111111",
		13440 => "11111111",
		13441 => "11111111",
		13442 => "11111111",
		13443 => "11111111",
		13444 => "11111111",
		13445 => "11111111",
		13446 => "11111111",
		13447 => "11111111",
		13448 => "11111111",
		13449 => "11111111",
		13450 => "11111111",
		13451 => "11111111",
		13452 => "11111111",
		13453 => "11111111",
		13454 => "11111111",
		13455 => "11111111",
		13456 => "11111111",
		13457 => "11111111",
		13458 => "11111111",
		13459 => "11111111",
		13460 => "11111111",
		13461 => "11111111",
		13462 => "11111111",
		13463 => "11111111",
		13464 => "11111111",
		13465 => "11111111",
		13466 => "11111111",
		13467 => "11111111",
		13468 => "11000101",
		13469 => "10000001",
		13470 => "10000111",
		13471 => "11101000",
		13472 => "11111111",
		13473 => "11111111",
		13474 => "11111111",
		13475 => "11111111",
		13476 => "11111111",
		13477 => "11111111",
		13478 => "11111111",
		13479 => "11111111",
		13480 => "11111111",
		13481 => "11111111",
		13482 => "11111111",
		13483 => "11111111",
		13484 => "11111111",
		13485 => "11011100",
		13486 => "01001101",
		13487 => "01111100",
		13488 => "11011100",
		13489 => "11111111",
		13490 => "11111111",
		13491 => "11111111",
		13492 => "11111111",
		13493 => "11111111",
		13494 => "11111111",
		13495 => "11111111",
		13496 => "11111111",
		13497 => "11111111",
		13498 => "11110011",
		13499 => "11001011",
		13500 => "10011000",
		13501 => "01100100",
		13502 => "01000111",
		13503 => "01000111",
		13504 => "01000111",
		13505 => "01000111",
		13506 => "01000111",
		13507 => "01100100",
		13508 => "10010011",
		13509 => "11000000",
		13510 => "11101110",
		13511 => "11111111",
		13512 => "11111111",
		13513 => "11111111",
		13514 => "11111111",
		13515 => "11111111",
		13516 => "11111111",
		13517 => "11111111",
		13518 => "11111111",
		13519 => "11110011",
		13520 => "10101110",
		13521 => "01010011",
		13522 => "01110101",
		13523 => "11111111",
		13524 => "11111111",
		13525 => "11111111",
		13526 => "11111111",
		13527 => "11111111",
		13528 => "11111111",
		13529 => "11111111",
		13530 => "11111111",
		13531 => "11111111",
		13532 => "11111111",
		13533 => "11111111",
		13534 => "11111111",
		13535 => "11111111",
		13536 => "11111111",
		13537 => "11111111",
		13538 => "10101110",
		13539 => "01000111",
		13540 => "01000111",
		13541 => "01000111",
		13542 => "01000111",
		13543 => "10101001",
		13544 => "11111111",
		13545 => "11111111",
		13546 => "11111111",
		13547 => "11111111",
		13548 => "11111111",
		13549 => "11111111",
		13550 => "11111111",
		13551 => "11111111",
		13552 => "11111111",
		13553 => "11111111",
		13554 => "11111111",
		13555 => "11111111",
		13556 => "11111111",
		13557 => "11111111",
		13558 => "11111111",
		13559 => "11111111",
		13560 => "11111111",
		13561 => "11111111",
		13562 => "11111111",
		13563 => "11111111",
		13564 => "11111111",
		13565 => "11111111",
		13566 => "11111111",
		13567 => "11111111",
		13568 => "11111111",
		13569 => "11111111",
		13570 => "11111111",
		13571 => "11111111",
		13572 => "11111111",
		13573 => "11111111",
		13574 => "11111111",
		13575 => "11111111",
		13576 => "11111111",
		13577 => "11111111",
		13578 => "11111111",
		13579 => "11111111",
		13580 => "11111111",
		13581 => "11111111",
		13582 => "11111111",
		13583 => "11111111",
		13584 => "11111111",
		13585 => "11111111",
		13586 => "11111111",
		13587 => "11111111",
		13588 => "11111111",
		13589 => "11111111",
		13590 => "11111111",
		13591 => "11111111",
		13592 => "11111111",
		13593 => "11111111",
		13594 => "11111111",
		13595 => "10111010",
		13596 => "01000111",
		13597 => "01000111",
		13598 => "01000111",
		13599 => "01011001",
		13600 => "11110011",
		13601 => "11111111",
		13602 => "11111111",
		13603 => "11111111",
		13604 => "11111111",
		13605 => "11111111",
		13606 => "11111111",
		13607 => "11111111",
		13608 => "11111111",
		13609 => "11111111",
		13610 => "11111111",
		13611 => "11111111",
		13612 => "11111111",
		13613 => "11111111",
		13614 => "10111010",
		13615 => "01011001",
		13616 => "01000111",
		13617 => "01011001",
		13618 => "01110101",
		13619 => "10010011",
		13620 => "10100011",
		13621 => "10100011",
		13622 => "10100011",
		13623 => "10100011",
		13624 => "01110101",
		13625 => "01011001",
		13626 => "01000111",
		13627 => "01000111",
		13628 => "01000111",
		13629 => "01110000",
		13630 => "10101001",
		13631 => "11011100",
		13632 => "11111111",
		13633 => "11011100",
		13634 => "10101110",
		13635 => "01111100",
		13636 => "01000111",
		13637 => "01000111",
		13638 => "01000111",
		13639 => "01000111",
		13640 => "01110101",
		13641 => "01111100",
		13642 => "10100011",
		13643 => "10100011",
		13644 => "10100011",
		13645 => "01110101",
		13646 => "01100100",
		13647 => "01000111",
		13648 => "01000111",
		13649 => "01110101",
		13650 => "11110011",
		13651 => "11111111",
		13652 => "11111111",
		13653 => "11111111",
		13654 => "11111111",
		13655 => "11111111",
		13656 => "11111111",
		13657 => "11111111",
		13658 => "11111111",
		13659 => "11111111",
		13660 => "11111111",
		13661 => "11111111",
		13662 => "11111111",
		13663 => "11111111",
		13664 => "11111111",
		13665 => "11111111",
		13666 => "10100011",
		13667 => "01000111",
		13668 => "01000111",
		13669 => "01000111",
		13670 => "01000111",
		13671 => "10010011",
		13672 => "11111111",
		13673 => "11111111",
		13674 => "11111111",
		13675 => "11111111",
		13676 => "11111111",
		13677 => "11111111",
		13678 => "11111111",
		13679 => "11111111",
		13680 => "11111111",
		13681 => "11111111",
		13682 => "11111111",
		13683 => "11111111",
		13684 => "11111111",
		13685 => "11111111",
		13686 => "11111111",
		13687 => "11111111",
		13688 => "11111111",
		13689 => "11111111",
		13690 => "11111111",
		13691 => "11111111",
		13692 => "11111111",
		13693 => "11111111",
		13694 => "11111111",
		13695 => "11111111",
		13696 => "11111111",
		13697 => "11111111",
		13698 => "11111111",
		13699 => "11111111",
		13700 => "11111111",
		13701 => "11111111",
		13702 => "11111111",
		13703 => "11111111",
		13704 => "11111111",
		13705 => "11111111",
		13706 => "11111111",
		13707 => "11111111",
		13708 => "11111111",
		13709 => "11111111",
		13710 => "11111111",
		13711 => "11111111",
		13712 => "11111111",
		13713 => "11111111",
		13714 => "11111111",
		13715 => "11111111",
		13716 => "11111111",
		13717 => "11111111",
		13718 => "11111111",
		13719 => "11111111",
		13720 => "11111111",
		13721 => "11111111",
		13722 => "11111111",
		13723 => "01110101",
		13724 => "01000111",
		13725 => "01000111",
		13726 => "01000111",
		13727 => "01000111",
		13728 => "11000000",
		13729 => "11111111",
		13730 => "11111111",
		13731 => "11111111",
		13732 => "11111111",
		13733 => "11111111",
		13734 => "11111111",
		13735 => "11111111",
		13736 => "11111111",
		13737 => "11111111",
		13738 => "11111111",
		13739 => "11111111",
		13740 => "11111111",
		13741 => "11111111",
		13742 => "11111111",
		13743 => "11110011",
		13744 => "10101001",
		13745 => "01111100",
		13746 => "01100100",
		13747 => "01000111",
		13748 => "01000111",
		13749 => "01000111",
		13750 => "01000111",
		13751 => "01000111",
		13752 => "01101010",
		13753 => "10000111",
		13754 => "10100011",
		13755 => "11010001",
		13756 => "11110011",
		13757 => "11111111",
		13758 => "11111111",
		13759 => "11111111",
		13760 => "11111111",
		13761 => "11111111",
		13762 => "11111111",
		13763 => "11111111",
		13764 => "11111001",
		13765 => "11010001",
		13766 => "10101110",
		13767 => "10100011",
		13768 => "01110101",
		13769 => "01101010",
		13770 => "01000111",
		13771 => "01000111",
		13772 => "01000111",
		13773 => "01110000",
		13774 => "10001100",
		13775 => "10100011",
		13776 => "11011100",
		13777 => "11111111",
		13778 => "11111111",
		13779 => "11111111",
		13780 => "11111111",
		13781 => "11111111",
		13782 => "11111111",
		13783 => "11111111",
		13784 => "11111111",
		13785 => "11111111",
		13786 => "11111111",
		13787 => "11111111",
		13788 => "11111111",
		13789 => "11111111",
		13790 => "11111111",
		13791 => "11111111",
		13792 => "11111111",
		13793 => "11111111",
		13794 => "11010111",
		13795 => "01000111",
		13796 => "01000111",
		13797 => "01000111",
		13798 => "01000111",
		13799 => "11011100",
		13800 => "11111111",
		13801 => "11111111",
		13802 => "11111111",
		13803 => "11111111",
		13804 => "11111111",
		13805 => "11111111",
		13806 => "11111111",
		13807 => "11111111",
		13808 => "11111111",
		13809 => "11111111",
		13810 => "11111111",
		13811 => "11111111",
		13812 => "11111111",
		13813 => "11111111",
		13814 => "11111111",
		13815 => "11111111",
		13816 => "11111111",
		13817 => "11111111",
		13818 => "11111111",
		13819 => "11111111",
		13820 => "11111111",
		13821 => "11111111",
		13822 => "11111111",
		13823 => "11111111",
		13824 => "11111111",
		13825 => "11111111",
		13826 => "11111111",
		13827 => "11111111",
		13828 => "11111111",
		13829 => "11111111",
		13830 => "11111111",
		13831 => "11111111",
		13832 => "11111111",
		13833 => "11111111",
		13834 => "11111111",
		13835 => "11111111",
		13836 => "11111111",
		13837 => "11111111",
		13838 => "11111111",
		13839 => "11111111",
		13840 => "11111111",
		13841 => "11111111",
		13842 => "11111111",
		13843 => "11111111",
		13844 => "11111111",
		13845 => "11111111",
		13846 => "11111111",
		13847 => "11111111",
		13848 => "11111111",
		13849 => "11111111",
		13850 => "11111111",
		13851 => "10011000",
		13852 => "01000111",
		13853 => "01000111",
		13854 => "01000111",
		13855 => "01000111",
		13856 => "11001011",
		13857 => "11111111",
		13858 => "11111111",
		13859 => "11111111",
		13860 => "11111111",
		13861 => "11111111",
		13862 => "11111111",
		13863 => "11111111",
		13864 => "11111111",
		13865 => "11111111",
		13866 => "11111111",
		13867 => "11111111",
		13868 => "11111111",
		13869 => "11111111",
		13870 => "11111111",
		13871 => "11111111",
		13872 => "11111111",
		13873 => "11111111",
		13874 => "11111111",
		13875 => "11111111",
		13876 => "11111111",
		13877 => "11111111",
		13878 => "11111111",
		13879 => "11111111",
		13880 => "11111111",
		13881 => "11111111",
		13882 => "11111111",
		13883 => "11111111",
		13884 => "11111111",
		13885 => "11111111",
		13886 => "11111111",
		13887 => "11111111",
		13888 => "11111111",
		13889 => "11111111",
		13890 => "11111111",
		13891 => "11111111",
		13892 => "11111111",
		13893 => "11111111",
		13894 => "11111111",
		13895 => "11111111",
		13896 => "11111111",
		13897 => "11111111",
		13898 => "11111111",
		13899 => "11111111",
		13900 => "11111111",
		13901 => "11111111",
		13902 => "11111111",
		13903 => "11111111",
		13904 => "11111111",
		13905 => "11111111",
		13906 => "11111111",
		13907 => "11111111",
		13908 => "11111111",
		13909 => "11111111",
		13910 => "11111111",
		13911 => "11111111",
		13912 => "11111111",
		13913 => "11111111",
		13914 => "11111111",
		13915 => "11111111",
		13916 => "11111111",
		13917 => "11111111",
		13918 => "11111111",
		13919 => "11111111",
		13920 => "11111111",
		13921 => "11111111",
		13922 => "11111111",
		13923 => "11011100",
		13924 => "10001100",
		13925 => "10000111",
		13926 => "11000101",
		13927 => "11111111",
		13928 => "11111111",
		13929 => "11111111",
		13930 => "11111111",
		13931 => "11111111",
		13932 => "11111111",
		13933 => "11111111",
		13934 => "11111111",
		13935 => "11111111",
		13936 => "11111111",
		13937 => "11111111",
		13938 => "11111111",
		13939 => "11111111",
		13940 => "11111111",
		13941 => "11111111",
		13942 => "11111111",
		13943 => "11111111",
		13944 => "11111111",
		13945 => "11111111",
		13946 => "11111111",
		13947 => "11111111",
		13948 => "11111111",
		13949 => "11111111",
		13950 => "11111111",
		13951 => "11111111",
		13952 => "11111111",
		13953 => "11111111",
		13954 => "11111111",
		13955 => "11111111",
		13956 => "11111111",
		13957 => "11111111",
		13958 => "11111111",
		13959 => "11111111",
		13960 => "11111111",
		13961 => "11111111",
		13962 => "11111111",
		13963 => "11111111",
		13964 => "11111111",
		13965 => "11111111",
		13966 => "11111111",
		13967 => "11111111",
		13968 => "11111111",
		13969 => "11111111",
		13970 => "11111111",
		13971 => "11111111",
		13972 => "11111111",
		13973 => "11111111",
		13974 => "11111111",
		13975 => "11111111",
		13976 => "11111111",
		13977 => "11111111",
		13978 => "11111111",
		13979 => "11101110",
		13980 => "01001101",
		13981 => "01000111",
		13982 => "01000111",
		13983 => "10010011",
		13984 => "11111111",
		13985 => "11111111",
		13986 => "11111111",
		13987 => "11111111",
		13988 => "11111111",
		13989 => "11111111",
		13990 => "11111111",
		13991 => "11111111",
		13992 => "11111111",
		13993 => "11111111",
		13994 => "11111111",
		13995 => "11111111",
		13996 => "11111111",
		13997 => "11111111",
		13998 => "11111111",
		13999 => "11111111",
		14000 => "11111111",
		14001 => "11111111",
		14002 => "11111111",
		14003 => "11111111",
		14004 => "11111111",
		14005 => "11111111",
		14006 => "11111111",
		14007 => "11111111",
		14008 => "11111111",
		14009 => "11111111",
		14010 => "11111111",
		14011 => "11111111",
		14012 => "11111111",
		14013 => "11111111",
		14014 => "11111111",
		14015 => "11111111",
		14016 => "11111111",
		14017 => "11111111",
		14018 => "11111111",
		14019 => "11111111",
		14020 => "11111111",
		14021 => "11111111",
		14022 => "11111111",
		14023 => "11111111",
		14024 => "11111111",
		14025 => "11111111",
		14026 => "11111111",
		14027 => "11111111",
		14028 => "11111111",
		14029 => "11111111",
		14030 => "11111111",
		14031 => "11111111",
		14032 => "11111111",
		14033 => "11111111",
		14034 => "11111111",
		14035 => "11111111",
		14036 => "11111111",
		14037 => "11111111",
		14038 => "11111111",
		14039 => "11111111",
		14040 => "11111111",
		14041 => "11111111",
		14042 => "11111111",
		14043 => "11111111",
		14044 => "11111111",
		14045 => "11111111",
		14046 => "11111111",
		14047 => "11111111",
		14048 => "11111111",
		14049 => "11111111",
		14050 => "11111111",
		14051 => "11111111",
		14052 => "11111111",
		14053 => "11111111",
		14054 => "11111111",
		14055 => "11111111",
		14056 => "11111111",
		14057 => "11111111",
		14058 => "11111111",
		14059 => "11111111",
		14060 => "11111111",
		14061 => "11111111",
		14062 => "11111111",
		14063 => "11111111",
		14064 => "11111111",
		14065 => "11111111",
		14066 => "11111111",
		14067 => "11111111",
		14068 => "11111111",
		14069 => "11111111",
		14070 => "11111111",
		14071 => "11111111",
		14072 => "11111111",
		14073 => "11111111",
		14074 => "11111111",
		14075 => "11111111",
		14076 => "11111111",
		14077 => "11111111",
		14078 => "11111111",
		14079 => "11111111",
		14080 => "11111111",
		14081 => "11111111",
		14082 => "11111111",
		14083 => "11111111",
		14084 => "11111111",
		14085 => "11111111",
		14086 => "11111111",
		14087 => "11111111",
		14088 => "11111111",
		14089 => "11111111",
		14090 => "11111111",
		14091 => "11111111",
		14092 => "11111111",
		14093 => "11111111",
		14094 => "11111111",
		14095 => "11111111",
		14096 => "11111111",
		14097 => "11111111",
		14098 => "11111111",
		14099 => "11111111",
		14100 => "11111111",
		14101 => "11111111",
		14102 => "11111111",
		14103 => "11111111",
		14104 => "11111111",
		14105 => "11111111",
		14106 => "11111111",
		14107 => "11111111",
		14108 => "11101110",
		14109 => "10111010",
		14110 => "11011100",
		14111 => "11111111",
		14112 => "11111111",
		14113 => "11111111",
		14114 => "11111111",
		14115 => "11111111",
		14116 => "11111111",
		14117 => "11111111",
		14118 => "11111111",
		14119 => "11111111",
		14120 => "11111111",
		14121 => "11111111",
		14122 => "11111111",
		14123 => "11111111",
		14124 => "11111111",
		14125 => "11111111",
		14126 => "11111111",
		14127 => "11111111",
		14128 => "11111111",
		14129 => "11111111",
		14130 => "11111111",
		14131 => "11111111",
		14132 => "11111111",
		14133 => "11111111",
		14134 => "11111111",
		14135 => "11111111",
		14136 => "11111111",
		14137 => "11111111",
		14138 => "11111111",
		14139 => "11111111",
		14140 => "11111111",
		14141 => "11111111",
		14142 => "11111111",
		14143 => "11111111",
		14144 => "11111111",
		14145 => "11111111",
		14146 => "11111111",
		14147 => "11111111",
		14148 => "11111111",
		14149 => "11111111",
		14150 => "11111111",
		14151 => "11111111",
		14152 => "11111111",
		14153 => "11111111",
		14154 => "11111111",
		14155 => "11111111",
		14156 => "11111111",
		14157 => "11111111",
		14158 => "11111111",
		14159 => "11111111",
		14160 => "11111111",
		14161 => "11111111",
		14162 => "11111111",
		14163 => "11111111",
		14164 => "11111111",
		14165 => "11111111",
		14166 => "11111111",
		14167 => "11111111",
		14168 => "11111111",
		14169 => "11111111",
		14170 => "11111111",
		14171 => "11111111",
		14172 => "11111111",
		14173 => "11111111",
		14174 => "11111111",
		14175 => "11111111",
		14176 => "11111111",
		14177 => "11111111",
		14178 => "11111111",
		14179 => "11111111",
		14180 => "11111111",
		14181 => "11111111",
		14182 => "11111111",
		14183 => "11111111",
		14184 => "11111111",
		14185 => "11111111",
		14186 => "11111111",
		14187 => "11111111",
		14188 => "11111111",
		14189 => "11111111",
		14190 => "11111111",
		14191 => "11111111",
		14192 => "11111111",
		14193 => "11111111",
		14194 => "11111111",
		14195 => "11111111",
		14196 => "11111111",
		14197 => "11111111",
		14198 => "11111111",
		14199 => "11111111",
		14200 => "11111111",
		14201 => "11111111",
		14202 => "11111111",
		14203 => "11111111",
		14204 => "11111111",
		14205 => "11111111",
		14206 => "11111111",
		14207 => "11111111",
		14208 => "11111111",
		14209 => "11111111",
		14210 => "11111111",
		14211 => "11111111",
		14212 => "11111111",
		14213 => "11111111",
		14214 => "11111111",
		14215 => "11111111",
		14216 => "11111111",
		14217 => "11111111",
		14218 => "11111111",
		14219 => "11111111",
		14220 => "11111111",
		14221 => "11111111",
		14222 => "11111111",
		14223 => "11111111",
		14224 => "11111111",
		14225 => "11111111",
		14226 => "11111111",
		14227 => "11111111",
		14228 => "11111111",
		14229 => "11111111",
		14230 => "11111111",
		14231 => "11111111",
		14232 => "11111111",
		14233 => "11111111",
		14234 => "11111111",
		14235 => "11111111",
		14236 => "11111111",
		14237 => "11111111",
		14238 => "11111111",
		14239 => "11111111",
		14240 => "11111111",
		14241 => "11111111",
		14242 => "11111111",
		14243 => "11111111",
		14244 => "11111111",
		14245 => "11111111",
		14246 => "11111111",
		14247 => "11111111",
		14248 => "11111111",
		14249 => "11111111",
		14250 => "11111111",
		14251 => "11111111",
		14252 => "11111111",
		14253 => "11111111",
		14254 => "11111111",
		14255 => "11111111",
		14256 => "11111111",
		14257 => "11111111",
		14258 => "11111111",
		14259 => "11111111",
		14260 => "11111111",
		14261 => "11111111",
		14262 => "11111111",
		14263 => "11111111",
		14264 => "11111111",
		14265 => "11111111",
		14266 => "11111111",
		14267 => "11111111",
		14268 => "11111111",
		14269 => "11111111",
		14270 => "11111111",
		14271 => "11111111",
		14272 => "11111111",
		14273 => "11111111",
		14274 => "11111111",
		14275 => "11111111",
		14276 => "11111111",
		14277 => "11111111",
		14278 => "11111111",
		14279 => "11111111",
		14280 => "11111111",
		14281 => "11111111",
		14282 => "11111111",
		14283 => "11111111",
		14284 => "11111111",
		14285 => "11111111",
		14286 => "11111111",
		14287 => "11111111",
		14288 => "11111111",
		14289 => "11111111",
		14290 => "11111111",
		14291 => "11111111",
		14292 => "11111111",
		14293 => "11111111",
		14294 => "11111111",
		14295 => "11111111",
		14296 => "11111111",
		14297 => "11111111",
		14298 => "11111111",
		14299 => "11111111",
		14300 => "11111111",
		14301 => "11111111",
		14302 => "11111111",
		14303 => "11111111",
		14304 => "11111111",
		14305 => "11111111",
		14306 => "11111111",
		14307 => "11111111",
		14308 => "11111111",
		14309 => "11111111",
		14310 => "11111111",
		14311 => "11111111",
		14312 => "11111111",
		14313 => "11111111",
		14314 => "11111111",
		14315 => "11111111",
		14316 => "11111111",
		14317 => "11111111",
		14318 => "11111111",
		14319 => "11111111",
		14320 => "11111111",
		14321 => "11111111",
		14322 => "11111111",
		14323 => "11111111",
		14324 => "11111111",
		14325 => "11111111",
		14326 => "11111111",
		14327 => "11111111",
		14328 => "11111111",
		14329 => "11111111",
		14330 => "11111111",
		14331 => "11111111",
		14332 => "11111111",
		14333 => "11111111",
		14334 => "11111111",
		14335 => "11111111",
		14336 => "11111111",
		14337 => "11111111",
		14338 => "11111111",
		14339 => "11111111",
		14340 => "11111111",
		14341 => "11111111",
		14342 => "11111111",
		14343 => "11111111",
		14344 => "11111111",
		14345 => "11111111",
		14346 => "11111111",
		14347 => "11111111",
		14348 => "11111111",
		14349 => "11111111",
		14350 => "11111111",
		14351 => "11111111",
		14352 => "11111111",
		14353 => "11111111",
		14354 => "11111111",
		14355 => "11111111",
		14356 => "11111111",
		14357 => "11111111",
		14358 => "11111111",
		14359 => "11111111",
		14360 => "11111111",
		14361 => "11111111",
		14362 => "11111111",
		14363 => "11111111",
		14364 => "11111111",
		14365 => "11111111",
		14366 => "11111111",
		14367 => "11111111",
		14368 => "11111111",
		14369 => "11111111",
		14370 => "11111111",
		14371 => "11111111",
		14372 => "11111111",
		14373 => "11111111",
		14374 => "11111111",
		14375 => "11111111",
		14376 => "11111111",
		14377 => "11111111",
		14378 => "11111111",
		14379 => "11111111",
		14380 => "11111111",
		14381 => "11111111",
		14382 => "11111111",
		14383 => "11111111",
		14384 => "11111111",
		14385 => "11111111",
		14386 => "11111111",
		14387 => "11111111",
		14388 => "11111111",
		14389 => "11111111",
		14390 => "11111111",
		14391 => "11111111",
		14392 => "11111111",
		14393 => "11111111",
		14394 => "11111111",
		14395 => "11111111",
		14396 => "11111111",
		14397 => "11111111",
		14398 => "11111111",
		14399 => "11111111",
		14400 => "11111111",
		14401 => "11111111",
		14402 => "11111111",
		14403 => "11111111",
		14404 => "11111111",
		14405 => "11111111",
		14406 => "11111111",
		14407 => "11111111",
		14408 => "11111111",
		14409 => "11111111",
		14410 => "11111111",
		14411 => "11111111",
		14412 => "11111111",
		14413 => "11111111",
		14414 => "11110011",
		14415 => "10111010",
		14416 => "10100011",
		14417 => "10100011",
		14418 => "11010001",
		14419 => "11111111",
		14420 => "11111111",
		14421 => "11111111",
		14422 => "11111111",
		14423 => "11111111",
		14424 => "11111111",
		14425 => "11111111",
		14426 => "11111111",
		14427 => "11111111",
		14428 => "11111111",
		14429 => "11111111",
		14430 => "11111111",
		14431 => "11111111",
		14432 => "11111111",
		14433 => "11111111",
		14434 => "11111111",
		14435 => "11111111",
		14436 => "11111111",
		14437 => "11111111",
		14438 => "11111111",
		14439 => "11111111",
		14440 => "11111111",
		14441 => "11111111",
		14442 => "11111111",
		14443 => "11111111",
		14444 => "11111111",
		14445 => "11111111",
		14446 => "11111111",
		14447 => "11111111",
		14448 => "11111111",
		14449 => "11111111",
		14450 => "11111111",
		14451 => "11111111",
		14452 => "11111111",
		14453 => "11111111",
		14454 => "11111111",
		14455 => "11111111",
		14456 => "11111111",
		14457 => "11111111",
		14458 => "11111111",
		14459 => "11111111",
		14460 => "11111111",
		14461 => "11111111",
		14462 => "11111111",
		14463 => "11111111",
		14464 => "11111111",
		14465 => "11111111",
		14466 => "11111111",
		14467 => "11111111",
		14468 => "11111111",
		14469 => "11111111",
		14470 => "11111111",
		14471 => "11111111",
		14472 => "11111111",
		14473 => "11111111",
		14474 => "11111111",
		14475 => "11111111",
		14476 => "11111111",
		14477 => "11111111",
		14478 => "11111111",
		14479 => "11111111",
		14480 => "11111111",
		14481 => "11111111",
		14482 => "11111111",
		14483 => "11111111",
		14484 => "11111111",
		14485 => "11111111",
		14486 => "11111111",
		14487 => "11111111",
		14488 => "11111111",
		14489 => "11111111",
		14490 => "11111111",
		14491 => "11111111",
		14492 => "11111111",
		14493 => "11111111",
		14494 => "11111111",
		14495 => "11111111",
		14496 => "11111111",
		14497 => "11111111",
		14498 => "11111111",
		14499 => "11111111",
		14500 => "11111111",
		14501 => "11111111",
		14502 => "11111111",
		14503 => "11111111",
		14504 => "11111111",
		14505 => "11111111",
		14506 => "11111111",
		14507 => "11111111",
		14508 => "11111111",
		14509 => "11011100",
		14510 => "10100011",
		14511 => "10100011",
		14512 => "10011000",
		14513 => "01110101",
		14514 => "01010011",
		14515 => "11111001",
		14516 => "11111111",
		14517 => "11111111",
		14518 => "11111111",
		14519 => "11111111",
		14520 => "11111111",
		14521 => "11111111",
		14522 => "11111111",
		14523 => "11111111",
		14524 => "11111111",
		14525 => "11111111",
		14526 => "11111111",
		14527 => "11111111",
		14528 => "11111111",
		14529 => "11111111",
		14530 => "11111111",
		14531 => "11111111",
		14532 => "11111111",
		14533 => "11111111",
		14534 => "11111111",
		14535 => "11111111",
		14536 => "11111111",
		14537 => "11111111",
		14538 => "11111111",
		14539 => "11111111",
		14540 => "11111001",
		14541 => "10100011",
		14542 => "01101010",
		14543 => "01110101",
		14544 => "01110101",
		14545 => "01000111",
		14546 => "01000111",
		14547 => "11010001",
		14548 => "11111111",
		14549 => "11111111",
		14550 => "11111111",
		14551 => "11111111",
		14552 => "11111111",
		14553 => "11111111",
		14554 => "11111111",
		14555 => "11111111",
		14556 => "11111111",
		14557 => "11111111",
		14558 => "11111111",
		14559 => "11111111",
		14560 => "11111111",
		14561 => "11111111",
		14562 => "11111111",
		14563 => "11111111",
		14564 => "11111111",
		14565 => "11111111",
		14566 => "11111111",
		14567 => "11111111",
		14568 => "11111111",
		14569 => "11111111",
		14570 => "11111111",
		14571 => "11111111",
		14572 => "11111111",
		14573 => "11111111",
		14574 => "11111111",
		14575 => "11111111",
		14576 => "11111111",
		14577 => "11111111",
		14578 => "11111111",
		14579 => "11111111",
		14580 => "11111111",
		14581 => "11111111",
		14582 => "11111111",
		14583 => "11111111",
		14584 => "11111111",
		14585 => "11111111",
		14586 => "11111111",
		14587 => "11111111",
		14588 => "11111111",
		14589 => "11111111",
		14590 => "11111111",
		14591 => "11111111",
		14592 => "11111111",
		14593 => "11111111",
		14594 => "11111111",
		14595 => "11111111",
		14596 => "11111111",
		14597 => "11111111",
		14598 => "11111111",
		14599 => "11111111",
		14600 => "11111111",
		14601 => "11111111",
		14602 => "11111111",
		14603 => "11111111",
		14604 => "11111111",
		14605 => "11111111",
		14606 => "11111111",
		14607 => "11111111",
		14608 => "11111111",
		14609 => "11111111",
		14610 => "11111111",
		14611 => "11111111",
		14612 => "11111111",
		14613 => "11111111",
		14614 => "11111111",
		14615 => "11111111",
		14616 => "11111111",
		14617 => "11111111",
		14618 => "11111111",
		14619 => "11111111",
		14620 => "11111111",
		14621 => "11111111",
		14622 => "11111111",
		14623 => "11111111",
		14624 => "11111111",
		14625 => "11111111",
		14626 => "11111111",
		14627 => "11111111",
		14628 => "11111111",
		14629 => "11111111",
		14630 => "11111111",
		14631 => "11111111",
		14632 => "11111111",
		14633 => "11111111",
		14634 => "11111111",
		14635 => "11111111",
		14636 => "11111111",
		14637 => "11101000",
		14638 => "11010001",
		14639 => "11000000",
		14640 => "10000111",
		14641 => "01000111",
		14642 => "10001100",
		14643 => "11111111",
		14644 => "11111111",
		14645 => "11111111",
		14646 => "11111111",
		14647 => "11111111",
		14648 => "11011100",
		14649 => "11010001",
		14650 => "11011100",
		14651 => "11111111",
		14652 => "11111111",
		14653 => "11111111",
		14654 => "11111111",
		14655 => "11111111",
		14656 => "11111111",
		14657 => "11111111",
		14658 => "11111111",
		14659 => "11111111",
		14660 => "11111111",
		14661 => "11111111",
		14662 => "11111111",
		14663 => "11100010",
		14664 => "11110011",
		14665 => "11111111",
		14666 => "11111111",
		14667 => "11111111",
		14668 => "10000001",
		14669 => "10000111",
		14670 => "11111111",
		14671 => "11111111",
		14672 => "11111111",
		14673 => "10011000",
		14674 => "01000111",
		14675 => "10000111",
		14676 => "11111111",
		14677 => "11111111",
		14678 => "11111111",
		14679 => "11111111",
		14680 => "11111111",
		14681 => "11111111",
		14682 => "11111111",
		14683 => "11111111",
		14684 => "11111111",
		14685 => "11111111",
		14686 => "11111111",
		14687 => "11111111",
		14688 => "11111111",
		14689 => "11111111",
		14690 => "11111111",
		14691 => "11111111",
		14692 => "11111111",
		14693 => "11111111",
		14694 => "11111111",
		14695 => "11111111",
		14696 => "11111111",
		14697 => "11111111",
		14698 => "11111111",
		14699 => "11111111",
		14700 => "11111111",
		14701 => "11111111",
		14702 => "11111111",
		14703 => "11111111",
		14704 => "11111111",
		14705 => "11111111",
		14706 => "11111111",
		14707 => "11111111",
		14708 => "11111111",
		14709 => "11111111",
		14710 => "11111111",
		14711 => "11111111",
		14712 => "11111111",
		14713 => "11111111",
		14714 => "11111111",
		14715 => "11111111",
		14716 => "11111111",
		14717 => "11111111",
		14718 => "11111111",
		14719 => "11111111",
		14720 => "11111111",
		14721 => "11111111",
		14722 => "11111111",
		14723 => "11111111",
		14724 => "11111111",
		14725 => "11111111",
		14726 => "11111111",
		14727 => "11111111",
		14728 => "11111111",
		14729 => "11111111",
		14730 => "11111111",
		14731 => "11111111",
		14732 => "11111111",
		14733 => "11111111",
		14734 => "11111111",
		14735 => "11111111",
		14736 => "11111111",
		14737 => "11111111",
		14738 => "11111111",
		14739 => "11111111",
		14740 => "11111111",
		14741 => "11111111",
		14742 => "11111111",
		14743 => "11111111",
		14744 => "11111111",
		14745 => "11111111",
		14746 => "11111111",
		14747 => "11111111",
		14748 => "11111111",
		14749 => "11111111",
		14750 => "11111111",
		14751 => "11111111",
		14752 => "11111111",
		14753 => "11111111",
		14754 => "11111111",
		14755 => "11111111",
		14756 => "11111111",
		14757 => "11111111",
		14758 => "11111111",
		14759 => "11111111",
		14760 => "11111111",
		14761 => "11111111",
		14762 => "11111111",
		14763 => "11111111",
		14764 => "11111111",
		14765 => "11111111",
		14766 => "11111111",
		14767 => "11111111",
		14768 => "01011001",
		14769 => "01011001",
		14770 => "11111001",
		14771 => "11111111",
		14772 => "11111111",
		14773 => "11111111",
		14774 => "11011100",
		14775 => "01101010",
		14776 => "11111111",
		14777 => "11111111",
		14778 => "11111111",
		14779 => "10011110",
		14780 => "01000111",
		14781 => "10100011",
		14782 => "11111111",
		14783 => "11111111",
		14784 => "11111111",
		14785 => "11111111",
		14786 => "11111111",
		14787 => "11111111",
		14788 => "11111111",
		14789 => "11111111",
		14790 => "10010011",
		14791 => "01000111",
		14792 => "10101110",
		14793 => "11111111",
		14794 => "11111111",
		14795 => "11111111",
		14796 => "11101000",
		14797 => "11000000",
		14798 => "11111111",
		14799 => "11111111",
		14800 => "11111111",
		14801 => "11011100",
		14802 => "01001101",
		14803 => "11101000",
		14804 => "11111111",
		14805 => "11111111",
		14806 => "11111111",
		14807 => "11111111",
		14808 => "11111111",
		14809 => "11111111",
		14810 => "11111111",
		14811 => "11111111",
		14812 => "11111111",
		14813 => "11111111",
		14814 => "11111111",
		14815 => "11111111",
		14816 => "11111111",
		14817 => "11111111",
		14818 => "11111111",
		14819 => "11111111",
		14820 => "11111111",
		14821 => "11111111",
		14822 => "11111111",
		14823 => "11111111",
		14824 => "11111111",
		14825 => "11111111",
		14826 => "11111111",
		14827 => "11111111",
		14828 => "11111111",
		14829 => "11111111",
		14830 => "11111111",
		14831 => "11111111",
		14832 => "11111111",
		14833 => "11111111",
		14834 => "11111111",
		14835 => "11111111",
		14836 => "11111111",
		14837 => "11111111",
		14838 => "11111111",
		14839 => "11111111",
		14840 => "11111111",
		14841 => "11111111",
		14842 => "11111111",
		14843 => "11111111",
		14844 => "11111111",
		14845 => "11111111",
		14846 => "11111111",
		14847 => "11111111",
		14848 => "11111111",
		14849 => "11111111",
		14850 => "11111111",
		14851 => "11111111",
		14852 => "11111111",
		14853 => "11111111",
		14854 => "11111111",
		14855 => "11111111",
		14856 => "11111111",
		14857 => "11111111",
		14858 => "11111111",
		14859 => "11111111",
		14860 => "11111111",
		14861 => "11111111",
		14862 => "11111111",
		14863 => "11111111",
		14864 => "11111111",
		14865 => "11111111",
		14866 => "11111111",
		14867 => "11111111",
		14868 => "11111111",
		14869 => "11111111",
		14870 => "11111111",
		14871 => "11111111",
		14872 => "11111111",
		14873 => "11111111",
		14874 => "11111111",
		14875 => "11111111",
		14876 => "11111111",
		14877 => "11111111",
		14878 => "11111111",
		14879 => "11111111",
		14880 => "11111111",
		14881 => "11111111",
		14882 => "11111111",
		14883 => "11111111",
		14884 => "11111111",
		14885 => "11111111",
		14886 => "11111111",
		14887 => "11111111",
		14888 => "11111111",
		14889 => "11111111",
		14890 => "11111111",
		14891 => "11111111",
		14892 => "11111111",
		14893 => "11111111",
		14894 => "11111111",
		14895 => "11010001",
		14896 => "01000111",
		14897 => "10010011",
		14898 => "11111111",
		14899 => "11111111",
		14900 => "11111111",
		14901 => "11111111",
		14902 => "11101000",
		14903 => "11010111",
		14904 => "11111111",
		14905 => "11111111",
		14906 => "11111111",
		14907 => "11010001",
		14908 => "01000111",
		14909 => "01110101",
		14910 => "11111111",
		14911 => "11111111",
		14912 => "11111111",
		14913 => "11111111",
		14914 => "11111111",
		14915 => "11111111",
		14916 => "11111111",
		14917 => "11010111",
		14918 => "01111100",
		14919 => "01000111",
		14920 => "10011000",
		14921 => "11111111",
		14922 => "11111111",
		14923 => "11111111",
		14924 => "11111111",
		14925 => "11111111",
		14926 => "11111111",
		14927 => "11111111",
		14928 => "11000101",
		14929 => "01100100",
		14930 => "10001100",
		14931 => "10101110",
		14932 => "11101110",
		14933 => "11111111",
		14934 => "11111111",
		14935 => "11111111",
		14936 => "11111111",
		14937 => "11111111",
		14938 => "11111111",
		14939 => "11111111",
		14940 => "11111111",
		14941 => "11111111",
		14942 => "11111111",
		14943 => "11111111",
		14944 => "11111111",
		14945 => "11111111",
		14946 => "11111111",
		14947 => "11111111",
		14948 => "11111111",
		14949 => "11111111",
		14950 => "11111111",
		14951 => "11111111",
		14952 => "11111111",
		14953 => "11111111",
		14954 => "11111111",
		14955 => "11111111",
		14956 => "11111111",
		14957 => "11111111",
		14958 => "11111111",
		14959 => "11111111",
		14960 => "11111111",
		14961 => "11111111",
		14962 => "11111111",
		14963 => "11111111",
		14964 => "11111111",
		14965 => "11111111",
		14966 => "11111111",
		14967 => "11111111",
		14968 => "11111111",
		14969 => "11111111",
		14970 => "11111111",
		14971 => "11111111",
		14972 => "11111111",
		14973 => "11111111",
		14974 => "11111111",
		14975 => "11111111",
		14976 => "11111111",
		14977 => "11111111",
		14978 => "11111111",
		14979 => "11111111",
		14980 => "11111111",
		14981 => "11111111",
		14982 => "11111111",
		14983 => "11111111",
		14984 => "11111111",
		14985 => "11111111",
		14986 => "11111111",
		14987 => "11111111",
		14988 => "11111111",
		14989 => "11111111",
		14990 => "11111111",
		14991 => "11111111",
		14992 => "11111111",
		14993 => "11111111",
		14994 => "11111111",
		14995 => "11111111",
		14996 => "11111111",
		14997 => "11111111",
		14998 => "11111111",
		14999 => "11111111",
		15000 => "11111111",
		15001 => "11111111",
		15002 => "11111111",
		15003 => "11111111",
		15004 => "11111111",
		15005 => "11111111",
		15006 => "11111111",
		15007 => "11111111",
		15008 => "11111111",
		15009 => "11111111",
		15010 => "11111111",
		15011 => "11111111",
		15012 => "11111111",
		15013 => "11111111",
		15014 => "11111111",
		15015 => "11111111",
		15016 => "11111111",
		15017 => "11111111",
		15018 => "11111111",
		15019 => "11111111",
		15020 => "11111111",
		15021 => "11111111",
		15022 => "11111111",
		15023 => "10010011",
		15024 => "01000111",
		15025 => "11010001",
		15026 => "11111111",
		15027 => "11111111",
		15028 => "11111111",
		15029 => "11111111",
		15030 => "11111111",
		15031 => "11111111",
		15032 => "11111111",
		15033 => "11111111",
		15034 => "11111111",
		15035 => "10101110",
		15036 => "01000111",
		15037 => "10001100",
		15038 => "11111111",
		15039 => "11111111",
		15040 => "11111111",
		15041 => "11111111",
		15042 => "11111111",
		15043 => "11111111",
		15044 => "11111001",
		15045 => "01110000",
		15046 => "11101000",
		15047 => "01011001",
		15048 => "10000111",
		15049 => "11111111",
		15050 => "11111111",
		15051 => "11111111",
		15052 => "11111111",
		15053 => "11111111",
		15054 => "11111111",
		15055 => "11111001",
		15056 => "10010011",
		15057 => "10100011",
		15058 => "10011000",
		15059 => "01000111",
		15060 => "01011110",
		15061 => "11101000",
		15062 => "11111111",
		15063 => "11111111",
		15064 => "11111111",
		15065 => "11111111",
		15066 => "11111111",
		15067 => "11111111",
		15068 => "11111111",
		15069 => "11111111",
		15070 => "11111111",
		15071 => "11111111",
		15072 => "11111111",
		15073 => "11111111",
		15074 => "11111111",
		15075 => "11111111",
		15076 => "11111111",
		15077 => "11111111",
		15078 => "11111111",
		15079 => "11111111",
		15080 => "11111111",
		15081 => "11111111",
		15082 => "11111111",
		15083 => "11111111",
		15084 => "11111111",
		15085 => "11111111",
		15086 => "11111111",
		15087 => "11111111",
		15088 => "11111111",
		15089 => "11111111",
		15090 => "11111111",
		15091 => "11111111",
		15092 => "11111111",
		15093 => "11111111",
		15094 => "11111111",
		15095 => "11111111",
		15096 => "11111111",
		15097 => "11111111",
		15098 => "11111111",
		15099 => "11111111",
		15100 => "11111111",
		15101 => "11111111",
		15102 => "11111111",
		15103 => "11111111",
		15104 => "11111111",
		15105 => "11111111",
		15106 => "11111111",
		15107 => "11111111",
		15108 => "11111111",
		15109 => "11111111",
		15110 => "11111111",
		15111 => "11111111",
		15112 => "11111111",
		15113 => "11111111",
		15114 => "11111111",
		15115 => "11111111",
		15116 => "11111111",
		15117 => "11111111",
		15118 => "11111111",
		15119 => "11111111",
		15120 => "11111111",
		15121 => "11111111",
		15122 => "11111111",
		15123 => "11111111",
		15124 => "11111111",
		15125 => "11111111",
		15126 => "11111111",
		15127 => "11111111",
		15128 => "11111111",
		15129 => "11111111",
		15130 => "11111111",
		15131 => "11111111",
		15132 => "11111111",
		15133 => "11111111",
		15134 => "11111111",
		15135 => "11111111",
		15136 => "11111111",
		15137 => "11111111",
		15138 => "11111111",
		15139 => "11111111",
		15140 => "11111111",
		15141 => "11111111",
		15142 => "11111111",
		15143 => "11111111",
		15144 => "11111111",
		15145 => "11111111",
		15146 => "11111111",
		15147 => "11111111",
		15148 => "11111111",
		15149 => "11111111",
		15150 => "11111111",
		15151 => "01011001",
		15152 => "01011001",
		15153 => "11111111",
		15154 => "11111111",
		15155 => "11111111",
		15156 => "11111111",
		15157 => "11111111",
		15158 => "11111111",
		15159 => "11111111",
		15160 => "11110011",
		15161 => "11010001",
		15162 => "11000000",
		15163 => "01011001",
		15164 => "01110101",
		15165 => "11101110",
		15166 => "11111111",
		15167 => "11111111",
		15168 => "11111111",
		15169 => "11111111",
		15170 => "11111111",
		15171 => "11111111",
		15172 => "10101001",
		15173 => "10011110",
		15174 => "11111111",
		15175 => "01110000",
		15176 => "01110101",
		15177 => "11111111",
		15178 => "11111111",
		15179 => "11111111",
		15180 => "11111111",
		15181 => "11111111",
		15182 => "11111111",
		15183 => "11111111",
		15184 => "11111111",
		15185 => "11111111",
		15186 => "11111111",
		15187 => "10101110",
		15188 => "01000111",
		15189 => "01101010",
		15190 => "11111111",
		15191 => "11111111",
		15192 => "11111111",
		15193 => "11111111",
		15194 => "11111111",
		15195 => "11111111",
		15196 => "11111111",
		15197 => "11111111",
		15198 => "11111111",
		15199 => "11111111",
		15200 => "11111111",
		15201 => "11111111",
		15202 => "11111111",
		15203 => "11111111",
		15204 => "11111111",
		15205 => "11111111",
		15206 => "11111111",
		15207 => "11111111",
		15208 => "11111111",
		15209 => "11111111",
		15210 => "11111111",
		15211 => "11111111",
		15212 => "11111111",
		15213 => "11111111",
		15214 => "11111111",
		15215 => "11111111",
		15216 => "11111111",
		15217 => "11111111",
		15218 => "11111111",
		15219 => "11111111",
		15220 => "11111111",
		15221 => "11111111",
		15222 => "11111111",
		15223 => "11111111",
		15224 => "11111111",
		15225 => "11111111",
		15226 => "11111111",
		15227 => "11111111",
		15228 => "11111111",
		15229 => "11111111",
		15230 => "11111111",
		15231 => "11111111",
		15232 => "11111111",
		15233 => "11111111",
		15234 => "11111111",
		15235 => "11111111",
		15236 => "11111111",
		15237 => "11111111",
		15238 => "11111111",
		15239 => "11111111",
		15240 => "11111111",
		15241 => "11111111",
		15242 => "11111111",
		15243 => "11111111",
		15244 => "11111111",
		15245 => "11111111",
		15246 => "11111111",
		15247 => "11111111",
		15248 => "11111111",
		15249 => "11111111",
		15250 => "11111111",
		15251 => "11111111",
		15252 => "11111111",
		15253 => "11111111",
		15254 => "11111111",
		15255 => "11111111",
		15256 => "11111111",
		15257 => "11111111",
		15258 => "11111111",
		15259 => "11111111",
		15260 => "11111111",
		15261 => "11111111",
		15262 => "11111111",
		15263 => "11111111",
		15264 => "11111111",
		15265 => "11111111",
		15266 => "11111111",
		15267 => "11111111",
		15268 => "11111111",
		15269 => "11111111",
		15270 => "11111111",
		15271 => "11111111",
		15272 => "11111111",
		15273 => "11111111",
		15274 => "11111111",
		15275 => "11111111",
		15276 => "11101110",
		15277 => "10001100",
		15278 => "01010011",
		15279 => "01000111",
		15280 => "01110000",
		15281 => "11111001",
		15282 => "11111111",
		15283 => "11111111",
		15284 => "11111111",
		15285 => "11111111",
		15286 => "11111111",
		15287 => "11111111",
		15288 => "11011100",
		15289 => "01100100",
		15290 => "01010011",
		15291 => "10101110",
		15292 => "11111111",
		15293 => "11111111",
		15294 => "11111111",
		15295 => "11111111",
		15296 => "11111111",
		15297 => "11111111",
		15298 => "11111111",
		15299 => "11101110",
		15300 => "01011110",
		15301 => "11111001",
		15302 => "11111111",
		15303 => "10000111",
		15304 => "01011110",
		15305 => "11111111",
		15306 => "11111111",
		15307 => "11111111",
		15308 => "11111111",
		15309 => "11111111",
		15310 => "11111111",
		15311 => "11111111",
		15312 => "11111111",
		15313 => "11111111",
		15314 => "11111111",
		15315 => "11111111",
		15316 => "01000111",
		15317 => "01011110",
		15318 => "11111111",
		15319 => "11111111",
		15320 => "11111111",
		15321 => "11111111",
		15322 => "11111111",
		15323 => "11111111",
		15324 => "11111111",
		15325 => "11111111",
		15326 => "11111111",
		15327 => "11111111",
		15328 => "11111111",
		15329 => "11111111",
		15330 => "11111111",
		15331 => "11111111",
		15332 => "11111111",
		15333 => "11111111",
		15334 => "11111111",
		15335 => "11111111",
		15336 => "11111111",
		15337 => "11111111",
		15338 => "11111111",
		15339 => "11111111",
		15340 => "11111111",
		15341 => "11111111",
		15342 => "11111111",
		15343 => "11111111",
		15344 => "11111111",
		15345 => "11111111",
		15346 => "11111111",
		15347 => "11111111",
		15348 => "11111111",
		15349 => "11111111",
		15350 => "11111111",
		15351 => "11111111",
		15352 => "11111111",
		15353 => "11111111",
		15354 => "11111111",
		15355 => "11111111",
		15356 => "11111111",
		15357 => "11111111",
		15358 => "11111111",
		15359 => "11111111",
		15360 => "11111111",
		15361 => "11111111",
		15362 => "11111111",
		15363 => "11111111",
		15364 => "11111111",
		15365 => "11111111",
		15366 => "11111111",
		15367 => "11111111",
		15368 => "11111111",
		15369 => "11111111",
		15370 => "11111111",
		15371 => "11111111",
		15372 => "11111111",
		15373 => "11111111",
		15374 => "11111111",
		15375 => "11111111",
		15376 => "11111111",
		15377 => "11111111",
		15378 => "11111111",
		15379 => "11111111",
		15380 => "11111111",
		15381 => "11111111",
		15382 => "11111111",
		15383 => "11111111",
		15384 => "11111111",
		15385 => "11111111",
		15386 => "11111111",
		15387 => "11111111",
		15388 => "11111111",
		15389 => "11111111",
		15390 => "11111111",
		15391 => "11111111",
		15392 => "11111111",
		15393 => "11111111",
		15394 => "11111111",
		15395 => "11111111",
		15396 => "11111111",
		15397 => "11111111",
		15398 => "11111111",
		15399 => "11111111",
		15400 => "11111111",
		15401 => "11111111",
		15402 => "11111111",
		15403 => "11111111",
		15404 => "11111111",
		15405 => "11111111",
		15406 => "11111111",
		15407 => "11001011",
		15408 => "10010011",
		15409 => "10000001",
		15410 => "11101110",
		15411 => "11111111",
		15412 => "11111111",
		15413 => "11111111",
		15414 => "11111111",
		15415 => "11111111",
		15416 => "11111111",
		15417 => "11111111",
		15418 => "11000101",
		15419 => "01011001",
		15420 => "10000001",
		15421 => "11111111",
		15422 => "11111111",
		15423 => "11111111",
		15424 => "11111111",
		15425 => "11111111",
		15426 => "11111111",
		15427 => "10000001",
		15428 => "10111010",
		15429 => "11111111",
		15430 => "11111111",
		15431 => "10011000",
		15432 => "01001101",
		15433 => "11111111",
		15434 => "11111111",
		15435 => "11111111",
		15436 => "11111111",
		15437 => "11111111",
		15438 => "11111111",
		15439 => "11111111",
		15440 => "11111111",
		15441 => "11111111",
		15442 => "11111111",
		15443 => "11101000",
		15444 => "01000111",
		15445 => "10011000",
		15446 => "11111111",
		15447 => "11111111",
		15448 => "11111111",
		15449 => "11111111",
		15450 => "11111111",
		15451 => "11111111",
		15452 => "11111111",
		15453 => "11111111",
		15454 => "11111111",
		15455 => "11111111",
		15456 => "11111111",
		15457 => "11111111",
		15458 => "11111111",
		15459 => "11111111",
		15460 => "11111111",
		15461 => "11111111",
		15462 => "11111111",
		15463 => "11111111",
		15464 => "11111111",
		15465 => "11111111",
		15466 => "11111111",
		15467 => "11111111",
		15468 => "11111111",
		15469 => "11111111",
		15470 => "11111111",
		15471 => "11111111",
		15472 => "11111111",
		15473 => "11111111",
		15474 => "11111111",
		15475 => "11111111",
		15476 => "11111111",
		15477 => "11111111",
		15478 => "11111111",
		15479 => "11111111",
		15480 => "11111111",
		15481 => "11111111",
		15482 => "11111111",
		15483 => "11111111",
		15484 => "11111111",
		15485 => "11111111",
		15486 => "11111111",
		15487 => "11111111",
		15488 => "11111111",
		15489 => "11111111",
		15490 => "11111111",
		15491 => "11111111",
		15492 => "11111111",
		15493 => "11111111",
		15494 => "11111111",
		15495 => "11111111",
		15496 => "11111111",
		15497 => "11111111",
		15498 => "11111111",
		15499 => "11111111",
		15500 => "11111111",
		15501 => "11111111",
		15502 => "11111111",
		15503 => "11111111",
		15504 => "11111111",
		15505 => "11111111",
		15506 => "11111111",
		15507 => "11111111",
		15508 => "11111111",
		15509 => "11111111",
		15510 => "11111111",
		15511 => "11111111",
		15512 => "11111111",
		15513 => "11111111",
		15514 => "11111111",
		15515 => "11111111",
		15516 => "11111111",
		15517 => "11111111",
		15518 => "11111111",
		15519 => "11111111",
		15520 => "11111111",
		15521 => "11111111",
		15522 => "11111111",
		15523 => "11111111",
		15524 => "11111111",
		15525 => "11111111",
		15526 => "11111111",
		15527 => "11111111",
		15528 => "11111111",
		15529 => "11111111",
		15530 => "11111111",
		15531 => "11111111",
		15532 => "11111111",
		15533 => "11111111",
		15534 => "11111111",
		15535 => "11111111",
		15536 => "11111111",
		15537 => "11111111",
		15538 => "11111111",
		15539 => "11111111",
		15540 => "11111111",
		15541 => "11111111",
		15542 => "11111111",
		15543 => "11111111",
		15544 => "11111111",
		15545 => "11111111",
		15546 => "11111111",
		15547 => "10001100",
		15548 => "01000111",
		15549 => "11000000",
		15550 => "11111111",
		15551 => "11111111",
		15552 => "11111111",
		15553 => "11111111",
		15554 => "11000101",
		15555 => "01111100",
		15556 => "11010111",
		15557 => "11010001",
		15558 => "10110100",
		15559 => "01110101",
		15560 => "01000111",
		15561 => "01110101",
		15562 => "11111111",
		15563 => "11111111",
		15564 => "11111111",
		15565 => "11111111",
		15566 => "11101000",
		15567 => "10000111",
		15568 => "11111111",
		15569 => "11111111",
		15570 => "11101110",
		15571 => "01101010",
		15572 => "01101010",
		15573 => "11110011",
		15574 => "11111111",
		15575 => "11111111",
		15576 => "11111111",
		15577 => "11111111",
		15578 => "11111111",
		15579 => "11111111",
		15580 => "11111111",
		15581 => "11111111",
		15582 => "11111111",
		15583 => "11111111",
		15584 => "11111111",
		15585 => "11111111",
		15586 => "11111111",
		15587 => "11111111",
		15588 => "11111111",
		15589 => "11111111",
		15590 => "11111111",
		15591 => "11111111",
		15592 => "11111111",
		15593 => "11111111",
		15594 => "11111111",
		15595 => "11111111",
		15596 => "11111111",
		15597 => "11111111",
		15598 => "11111111",
		15599 => "11111111",
		15600 => "11111111",
		15601 => "11111111",
		15602 => "11111111",
		15603 => "11111111",
		15604 => "11111111",
		15605 => "11111111",
		15606 => "11111111",
		15607 => "11111111",
		15608 => "11111111",
		15609 => "11111111",
		15610 => "11111111",
		15611 => "11111111",
		15612 => "11111111",
		15613 => "11111111",
		15614 => "11111111",
		15615 => "11111111",
		15616 => "11111111",
		15617 => "11111111",
		15618 => "11111111",
		15619 => "11111111",
		15620 => "11111111",
		15621 => "11111111",
		15622 => "11111111",
		15623 => "11111111",
		15624 => "11111111",
		15625 => "11111111",
		15626 => "11111111",
		15627 => "11111111",
		15628 => "11111111",
		15629 => "11111111",
		15630 => "11111111",
		15631 => "11111111",
		15632 => "11111111",
		15633 => "11111111",
		15634 => "11111111",
		15635 => "11111111",
		15636 => "11111111",
		15637 => "11111111",
		15638 => "11111111",
		15639 => "11111111",
		15640 => "11111111",
		15641 => "11111111",
		15642 => "11111111",
		15643 => "11111111",
		15644 => "11111111",
		15645 => "11111111",
		15646 => "11111111",
		15647 => "11111111",
		15648 => "11111111",
		15649 => "11111111",
		15650 => "11111111",
		15651 => "11111111",
		15652 => "11111111",
		15653 => "11111111",
		15654 => "11111111",
		15655 => "11111111",
		15656 => "11111111",
		15657 => "11111111",
		15658 => "11111111",
		15659 => "11111111",
		15660 => "11111111",
		15661 => "11111111",
		15662 => "11111111",
		15663 => "11111111",
		15664 => "11111111",
		15665 => "11111111",
		15666 => "11111111",
		15667 => "11111111",
		15668 => "11111111",
		15669 => "11111111",
		15670 => "10110100",
		15671 => "11111111",
		15672 => "11111111",
		15673 => "11111111",
		15674 => "11111111",
		15675 => "10011110",
		15676 => "01000111",
		15677 => "10101001",
		15678 => "11111111",
		15679 => "11111111",
		15680 => "11111111",
		15681 => "11111111",
		15682 => "01011001",
		15683 => "01000111",
		15684 => "01000111",
		15685 => "01010011",
		15686 => "01110101",
		15687 => "01101010",
		15688 => "01000111",
		15689 => "10001100",
		15690 => "11111111",
		15691 => "11111111",
		15692 => "11111111",
		15693 => "11111111",
		15694 => "11111111",
		15695 => "01011110",
		15696 => "10000111",
		15697 => "10000001",
		15698 => "01011001",
		15699 => "10101110",
		15700 => "11111001",
		15701 => "11111111",
		15702 => "11111111",
		15703 => "11111111",
		15704 => "11111111",
		15705 => "11111111",
		15706 => "11111111",
		15707 => "11111111",
		15708 => "11111111",
		15709 => "11111111",
		15710 => "11111111",
		15711 => "11111111",
		15712 => "11111111",
		15713 => "11111111",
		15714 => "11111111",
		15715 => "11111111",
		15716 => "11111111",
		15717 => "11111111",
		15718 => "11111111",
		15719 => "11111111",
		15720 => "11111111",
		15721 => "11111111",
		15722 => "11111111",
		15723 => "11111111",
		15724 => "11111111",
		15725 => "11111111",
		15726 => "11111111",
		15727 => "11111111",
		15728 => "11111111",
		15729 => "11111111",
		15730 => "11111111",
		15731 => "11111111",
		15732 => "11111111",
		15733 => "11111111",
		15734 => "11111111",
		15735 => "11111111",
		15736 => "11111111",
		15737 => "11111111",
		15738 => "11111111",
		15739 => "11111111",
		15740 => "11111111",
		15741 => "11111111",
		15742 => "11111111",
		15743 => "11111111",
		15744 => "11111111",
		15745 => "11111111",
		15746 => "11111111",
		15747 => "11111111",
		15748 => "11111111",
		15749 => "11111111",
		15750 => "11111111",
		15751 => "11111111",
		15752 => "11111111",
		15753 => "11111111",
		15754 => "11111111",
		15755 => "11111111",
		15756 => "11111111",
		15757 => "11111111",
		15758 => "11111111",
		15759 => "11111111",
		15760 => "11111111",
		15761 => "11111111",
		15762 => "11111111",
		15763 => "11111111",
		15764 => "11111111",
		15765 => "11111111",
		15766 => "11111111",
		15767 => "11111111",
		15768 => "11111111",
		15769 => "11111111",
		15770 => "11111111",
		15771 => "11111111",
		15772 => "11111111",
		15773 => "11111111",
		15774 => "11111111",
		15775 => "11111111",
		15776 => "11111111",
		15777 => "11111111",
		15778 => "11111111",
		15779 => "11111111",
		15780 => "11111111",
		15781 => "11111111",
		15782 => "11111111",
		15783 => "11111111",
		15784 => "11111111",
		15785 => "11111111",
		15786 => "11111111",
		15787 => "11111111",
		15788 => "11111111",
		15789 => "11111111",
		15790 => "11111111",
		15791 => "11111111",
		15792 => "11111111",
		15793 => "11111111",
		15794 => "11111111",
		15795 => "11111111",
		15796 => "11111111",
		15797 => "11111111",
		15798 => "01110101",
		15799 => "11111111",
		15800 => "11111111",
		15801 => "11111111",
		15802 => "11100010",
		15803 => "01001101",
		15804 => "01000111",
		15805 => "11100010",
		15806 => "11111111",
		15807 => "11111111",
		15808 => "11111111",
		15809 => "11111111",
		15810 => "11010001",
		15811 => "11110011",
		15812 => "11111111",
		15813 => "11111111",
		15814 => "11111111",
		15815 => "11010001",
		15816 => "01000111",
		15817 => "11000101",
		15818 => "11111111",
		15819 => "11111111",
		15820 => "11111111",
		15821 => "11111111",
		15822 => "11111111",
		15823 => "11000000",
		15824 => "10101001",
		15825 => "11011100",
		15826 => "11111111",
		15827 => "11111111",
		15828 => "11111111",
		15829 => "11111111",
		15830 => "11111111",
		15831 => "11111111",
		15832 => "11111111",
		15833 => "11111111",
		15834 => "11111111",
		15835 => "11111111",
		15836 => "11111111",
		15837 => "11111111",
		15838 => "11111111",
		15839 => "11111111",
		15840 => "11111111",
		15841 => "11111111",
		15842 => "11111111",
		15843 => "11111111",
		15844 => "11111111",
		15845 => "11111111",
		15846 => "11111111",
		15847 => "11111111",
		15848 => "11111111",
		15849 => "11111111",
		15850 => "11111111",
		15851 => "11111111",
		15852 => "11111111",
		15853 => "11111111",
		15854 => "11111111",
		15855 => "11111111",
		15856 => "11111111",
		15857 => "11111111",
		15858 => "11111111",
		15859 => "11111111",
		15860 => "11111111",
		15861 => "11111111",
		15862 => "11111111",
		15863 => "11111111",
		15864 => "11111111",
		15865 => "11111111",
		15866 => "11111111",
		15867 => "11111111",
		15868 => "11111111",
		15869 => "11111111",
		15870 => "11111111",
		15871 => "11111111",
		15872 => "11111111",
		15873 => "11111111",
		15874 => "11111111",
		15875 => "11111111",
		15876 => "11111111",
		15877 => "11111111",
		15878 => "11111111",
		15879 => "11111111",
		15880 => "11111111",
		15881 => "11111111",
		15882 => "11111111",
		15883 => "11111111",
		15884 => "11111111",
		15885 => "11111111",
		15886 => "11111111",
		15887 => "11111111",
		15888 => "11111111",
		15889 => "11111111",
		15890 => "11111111",
		15891 => "11111111",
		15892 => "11111111",
		15893 => "11111111",
		15894 => "11111111",
		15895 => "11111111",
		15896 => "11111111",
		15897 => "11111111",
		15898 => "11111111",
		15899 => "11111111",
		15900 => "11111111",
		15901 => "11111111",
		15902 => "11111111",
		15903 => "11111111",
		15904 => "11111111",
		15905 => "11111111",
		15906 => "11111111",
		15907 => "11111111",
		15908 => "11111111",
		15909 => "11111111",
		15910 => "11111111",
		15911 => "11111111",
		15912 => "11111111",
		15913 => "11111111",
		15914 => "11111111",
		15915 => "11111111",
		15916 => "11111111",
		15917 => "11111111",
		15918 => "11111111",
		15919 => "11111111",
		15920 => "11111111",
		15921 => "11111111",
		15922 => "11111111",
		15923 => "11111111",
		15924 => "11111111",
		15925 => "11111111",
		15926 => "01001101",
		15927 => "10000001",
		15928 => "10100011",
		15929 => "10010011",
		15930 => "01011001",
		15931 => "01010011",
		15932 => "11000101",
		15933 => "11111111",
		15934 => "11111111",
		15935 => "11111111",
		15936 => "11111111",
		15937 => "11111111",
		15938 => "11111111",
		15939 => "11111111",
		15940 => "11111111",
		15941 => "11111111",
		15942 => "11111111",
		15943 => "11101000",
		15944 => "01000111",
		15945 => "10110100",
		15946 => "11111111",
		15947 => "11111111",
		15948 => "11111111",
		15949 => "11111111",
		15950 => "11111111",
		15951 => "11111111",
		15952 => "11111111",
		15953 => "11111111",
		15954 => "11111111",
		15955 => "11111111",
		15956 => "11111111",
		15957 => "11111111",
		15958 => "11111111",
		15959 => "11111111",
		15960 => "11111111",
		15961 => "11111111",
		15962 => "11111111",
		15963 => "11111111",
		15964 => "11111111",
		15965 => "11111111",
		15966 => "11111111",
		15967 => "11111111",
		15968 => "11111111",
		15969 => "11111111",
		15970 => "11111111",
		15971 => "11111111",
		15972 => "11111111",
		15973 => "11111111",
		15974 => "11111111",
		15975 => "11111111",
		15976 => "11111111",
		15977 => "11111111",
		15978 => "11111111",
		15979 => "11111111",
		15980 => "11111111",
		15981 => "11111111",
		15982 => "11111111",
		15983 => "11111111",
		15984 => "11111111",
		15985 => "11111111",
		15986 => "11111111",
		15987 => "11111111",
		15988 => "11111111",
		15989 => "11111111",
		15990 => "11111111",
		15991 => "11111111",
		15992 => "11111111",
		15993 => "11111111",
		15994 => "11111111",
		15995 => "11111111",
		15996 => "11111111",
		15997 => "11111111",
		15998 => "11111111",
		15999 => "11111111",
		16000 => "11111111",
		16001 => "11111111",
		16002 => "11111111",
		16003 => "11111111",
		16004 => "11111111",
		16005 => "11111111",
		16006 => "11111111",
		16007 => "11111111",
		16008 => "11111111",
		16009 => "11111111",
		16010 => "11111111",
		16011 => "11111111",
		16012 => "11111111",
		16013 => "11111111",
		16014 => "11111111",
		16015 => "11111111",
		16016 => "11111111",
		16017 => "11111111",
		16018 => "11111111",
		16019 => "11111111",
		16020 => "11111111",
		16021 => "11111111",
		16022 => "11111111",
		16023 => "11111111",
		16024 => "11111111",
		16025 => "11111111",
		16026 => "11111111",
		16027 => "11111111",
		16028 => "11111111",
		16029 => "11111111",
		16030 => "11111111",
		16031 => "11111111",
		16032 => "11111111",
		16033 => "11111111",
		16034 => "11111111",
		16035 => "11111111",
		16036 => "11111111",
		16037 => "11111111",
		16038 => "11111111",
		16039 => "11111111",
		16040 => "11111111",
		16041 => "11111111",
		16042 => "11111111",
		16043 => "11111111",
		16044 => "11111111",
		16045 => "11111111",
		16046 => "11111111",
		16047 => "11111111",
		16048 => "11111111",
		16049 => "11111111",
		16050 => "11111111",
		16051 => "11111111",
		16052 => "11111111",
		16053 => "11111111",
		16054 => "11111111",
		16055 => "11111111",
		16056 => "11111111",
		16057 => "11111111",
		16058 => "11111111",
		16059 => "11111111",
		16060 => "11111111",
		16061 => "11111111",
		16062 => "11111111",
		16063 => "11111111",
		16064 => "11111111",
		16065 => "11111111",
		16066 => "11111111",
		16067 => "11111111",
		16068 => "11111111",
		16069 => "11111111",
		16070 => "11111111",
		16071 => "11111111",
		16072 => "11111111",
		16073 => "11111111",
		16074 => "11111111",
		16075 => "11111111",
		16076 => "11111111",
		16077 => "11111111",
		16078 => "11111111",
		16079 => "11111111",
		16080 => "11111111",
		16081 => "11111111",
		16082 => "11111111",
		16083 => "11111111",
		16084 => "11111111",
		16085 => "11111111",
		16086 => "11111111",
		16087 => "11111111",
		16088 => "11111111",
		16089 => "11111111",
		16090 => "11111111",
		16091 => "11111111",
		16092 => "11111111",
		16093 => "11111111",
		16094 => "11111111",
		16095 => "11111111",
		16096 => "11111111",
		16097 => "11111111",
		16098 => "11111111",
		16099 => "11111111",
		16100 => "11111111",
		16101 => "11111111",
		16102 => "11111111",
		16103 => "11111111",
		16104 => "11111111",
		16105 => "11111111",
		16106 => "11111111",
		16107 => "11111111",
		16108 => "11111111",
		16109 => "11111111",
		16110 => "11111111",
		16111 => "11111111",
		16112 => "11111111",
		16113 => "11111111",
		16114 => "11111111",
		16115 => "11111111",
		16116 => "11111111",
		16117 => "11111111",
		16118 => "11111111",
		16119 => "11111111",
		16120 => "11111111",
		16121 => "11111111",
		16122 => "11111111",
		16123 => "11111111",
		16124 => "11111111",
		16125 => "11111111",
		16126 => "11111111",
		16127 => "11111111",
		16128 => "11111111",
		16129 => "11111111",
		16130 => "11111111",
		16131 => "11111111",
		16132 => "11111111",
		16133 => "11111111",
		16134 => "11111111",
		16135 => "11111111",
		16136 => "11111111",
		16137 => "11111111",
		16138 => "11111111",
		16139 => "11111111",
		16140 => "11111111",
		16141 => "11111111",
		16142 => "11111111",
		16143 => "11111111",
		16144 => "11111111",
		16145 => "11111111",
		16146 => "11111111",
		16147 => "11111111",
		16148 => "11111111",
		16149 => "11111111",
		16150 => "11111111",
		16151 => "11111111",
		16152 => "11111111",
		16153 => "11111111",
		16154 => "11111111",
		16155 => "11111111",
		16156 => "11111111",
		16157 => "11111111",
		16158 => "11111111",
		16159 => "11111111",
		16160 => "11111111",
		16161 => "11111111",
		16162 => "11111111",
		16163 => "11111111",
		16164 => "11111111",
		16165 => "11111111",
		16166 => "11111111",
		16167 => "11111111",
		16168 => "11111111",
		16169 => "11111111",
		16170 => "11111111",
		16171 => "11111111",
		16172 => "11111111",
		16173 => "11111111",
		16174 => "11111111",
		16175 => "11111111",
		16176 => "11111111",
		16177 => "11111111",
		16178 => "11111111",
		16179 => "11111111",
		16180 => "11111111",
		16181 => "11111111",
		16182 => "11111111",
		16183 => "11111111",
		16184 => "11111111",
		16185 => "11111111",
		16186 => "11111111",
		16187 => "11111111",
		16188 => "11111111",
		16189 => "11111111",
		16190 => "11111111",
		16191 => "11111111",
		16192 => "11111111",
		16193 => "11111111",
		16194 => "11111111",
		16195 => "11111111",
		16196 => "11111111",
		16197 => "11111111",
		16198 => "11111111",
		16199 => "11111111",
		16200 => "11111111",
		16201 => "11111111",
		16202 => "11111111",
		16203 => "11111111",
		16204 => "11111111",
		16205 => "11111111",
		16206 => "11111111",
		16207 => "11111111",
		16208 => "11111111",
		16209 => "11111111",
		16210 => "11111111",
		16211 => "11111111",
		16212 => "11111111",
		16213 => "11111111",
		16214 => "11111111",
		16215 => "11111111",
		16216 => "11111111",
		16217 => "11111111",
		16218 => "11111111",
		16219 => "11111111",
		16220 => "11111111",
		16221 => "11111111",
		16222 => "11111111",
		16223 => "11111111",
		16224 => "11111111",
		16225 => "11111111",
		16226 => "11111111",
		16227 => "11111111",
		16228 => "11111111",
		16229 => "11111111",
		16230 => "11111111",
		16231 => "11111111",
		16232 => "11111111",
		16233 => "11111111",
		16234 => "11111111",
		16235 => "11111111",
		16236 => "11111111",
		16237 => "11111111",
		16238 => "11111111",
		16239 => "11111111",
		16240 => "11111111",
		16241 => "11111111",
		16242 => "11111111",
		16243 => "11111111",
		16244 => "11111111",
		16245 => "11111111",
		16246 => "11111111",
		16247 => "11111111",
		16248 => "11111111",
		16249 => "11111111",
		16250 => "11111111",
		16251 => "11111111",
		16252 => "11111111",
		16253 => "11111111",
		16254 => "11111111",
		16255 => "11111111",
		16256 => "11111111",
		16257 => "11111111",
		16258 => "11111111",
		16259 => "11111111",
		16260 => "11111111",
		16261 => "11111111",
		16262 => "11111111",
		16263 => "11111111",
		16264 => "11111111",
		16265 => "11111111",
		16266 => "11111111",
		16267 => "11111111",
		16268 => "11111111",
		16269 => "11111111",
		16270 => "11111111",
		16271 => "11111111",
		16272 => "11111111",
		16273 => "11111111",
		16274 => "11111111",
		16275 => "11111111",
		16276 => "11111111",
		16277 => "11111111",
		16278 => "11111111",
		16279 => "11111111",
		16280 => "11111111",
		16281 => "11111111",
		16282 => "11111111",
		16283 => "11111111",
		16284 => "11111111",
		16285 => "11111111",
		16286 => "11111111",
		16287 => "11111111",
		16288 => "11111111",
		16289 => "11111111",
		16290 => "11111111",
		16291 => "11111111",
		16292 => "11111111",
		16293 => "11111111",
		16294 => "11111111",
		16295 => "11111111",
		16296 => "11111111",
		16297 => "11111111",
		16298 => "11111111",
		16299 => "11111111",
		16300 => "11111111",
		16301 => "11111111",
		16302 => "11111111",
		16303 => "11111111",
		16304 => "11111111",
		16305 => "11111111",
		16306 => "11111111",
		16307 => "11111111",
		16308 => "11111111",
		16309 => "11111111",
		16310 => "11111111",
		16311 => "11111111",
		16312 => "11111111",
		16313 => "11111111",
		16314 => "11111111",
		16315 => "11111111",
		16316 => "11111111",
		16317 => "11111111",
		16318 => "11111111",
		16319 => "11111111",
		16320 => "11111111",
		16321 => "11111111",
		16322 => "11111111",
		16323 => "11111111",
		16324 => "11111111",
		16325 => "11111111",
		16326 => "11111111",
		16327 => "11111111",
		16328 => "11111111",
		16329 => "11111111",
		16330 => "11111111",
		16331 => "11111111",
		16332 => "11111111",
		16333 => "11111111",
		16334 => "11111111",
		16335 => "11111111",
		16336 => "11111111",
		16337 => "11111111",
		16338 => "11111111",
		16339 => "11111111",
		16340 => "11111111",
		16341 => "11111111",
		16342 => "11111111",
		16343 => "11111111",
		16344 => "11111111",
		16345 => "11111111",
		16346 => "11111111",
		16347 => "11111111",
		16348 => "11111111",
		16349 => "11111111",
		16350 => "11111111",
		16351 => "11111111",
		16352 => "11111111",
		16353 => "11111111",
		16354 => "11111111",
		16355 => "11111111",
		16356 => "11111111",
		16357 => "11111111",
		16358 => "11111111",
		16359 => "11111111",
		16360 => "11111111",
		16361 => "11111111",
		16362 => "11111111",
		16363 => "11111111",
		16364 => "11111111",
		16365 => "11111111",
		16366 => "11111111",
		16367 => "11111111",
		16368 => "11111111",
		16369 => "11111111",
		16370 => "11111111",
		16371 => "11111111",
		16372 => "11111111",
		16373 => "11111111",
		16374 => "11111111",
		16375 => "11111111",
		16376 => "11111111",
		16377 => "11111111",
		16378 => "11111111",
		16379 => "11111111",
		16380 => "11111111",
		16381 => "11111111",
		16382 => "11111111",
		16383 => "11111111"
	);

begin

	value <= ROM( to_integer( unsigned(address) ) );

end architecture;
