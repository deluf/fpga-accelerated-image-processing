
library IEEE;
	use IEEE.std_logic_1164.all;
	use IEEE.numeric_std.all;

entity Wrapper_SmallROM_SmallPixels is
	port (
		address	: in	std_logic_vector(7 downto 0);
		value	: out	std_logic_vector(3 downto 0)
	);
end entity;

architecture Arch of Wrapper_SmallROM_SmallPixels is

	type ROM_t is array (natural range 0 to 255) of std_logic_vector(3 downto 0);
	constant ROM: ROM_t := (
		0 => "1111",
		1 => "1111",
		2 => "1111",
		3 => "1111",
		4 => "1111",
		5 => "1111",
		6 => "1111",
		7 => "1111",
		8 => "1111",
		9 => "1111",
		10 => "1111",
		11 => "1111",
		12 => "1111",
		13 => "1111",
		14 => "1111",
		15 => "1111",
		16 => "1110",
		17 => "1110",
		18 => "1110",
		19 => "1110",
		20 => "1110",
		21 => "1110",
		22 => "1110",
		23 => "1110",
		24 => "1110",
		25 => "1110",
		26 => "1110",
		27 => "1110",
		28 => "1110",
		29 => "1110",
		30 => "1110",
		31 => "1110",
		32 => "1101",
		33 => "1101",
		34 => "1101",
		35 => "1101",
		36 => "1101",
		37 => "1101",
		38 => "1101",
		39 => "1101",
		40 => "1101",
		41 => "1101",
		42 => "1101",
		43 => "1101",
		44 => "1101",
		45 => "1101",
		46 => "1101",
		47 => "1101",
		48 => "1100",
		49 => "1100",
		50 => "1100",
		51 => "1100",
		52 => "1100",
		53 => "1100",
		54 => "1100",
		55 => "1100",
		56 => "1100",
		57 => "1100",
		58 => "1100",
		59 => "1100",
		60 => "1100",
		61 => "1100",
		62 => "1100",
		63 => "1100",
		64 => "1011",
		65 => "1011",
		66 => "1011",
		67 => "1011",
		68 => "1011",
		69 => "1011",
		70 => "1011",
		71 => "1011",
		72 => "1011",
		73 => "1011",
		74 => "1011",
		75 => "1011",
		76 => "1011",
		77 => "1011",
		78 => "1011",
		79 => "1011",
		80 => "1010",
		81 => "1010",
		82 => "1010",
		83 => "1010",
		84 => "1010",
		85 => "1010",
		86 => "1010",
		87 => "1010",
		88 => "1010",
		89 => "1010",
		90 => "1010",
		91 => "1010",
		92 => "1010",
		93 => "1010",
		94 => "1010",
		95 => "1010",
		96 => "1001",
		97 => "1001",
		98 => "1001",
		99 => "1001",
		100 => "1001",
		101 => "1001",
		102 => "1001",
		103 => "1001",
		104 => "1001",
		105 => "1001",
		106 => "1001",
		107 => "1001",
		108 => "1001",
		109 => "1001",
		110 => "1001",
		111 => "1001",
		112 => "1000",
		113 => "1000",
		114 => "1000",
		115 => "1000",
		116 => "1000",
		117 => "1000",
		118 => "1000",
		119 => "1000",
		120 => "1000",
		121 => "1000",
		122 => "1000",
		123 => "1000",
		124 => "1000",
		125 => "1000",
		126 => "1000",
		127 => "1000",
		128 => "0111",
		129 => "0111",
		130 => "0111",
		131 => "0111",
		132 => "0111",
		133 => "0111",
		134 => "0111",
		135 => "0111",
		136 => "0111",
		137 => "0111",
		138 => "0111",
		139 => "0111",
		140 => "0111",
		141 => "0111",
		142 => "0111",
		143 => "0111",
		144 => "0110",
		145 => "0110",
		146 => "0110",
		147 => "0110",
		148 => "0110",
		149 => "0110",
		150 => "0110",
		151 => "0110",
		152 => "0110",
		153 => "0110",
		154 => "0110",
		155 => "0110",
		156 => "0110",
		157 => "0110",
		158 => "0110",
		159 => "0110",
		160 => "0101",
		161 => "0101",
		162 => "0101",
		163 => "0101",
		164 => "0101",
		165 => "0101",
		166 => "0101",
		167 => "0101",
		168 => "0101",
		169 => "0101",
		170 => "0101",
		171 => "0101",
		172 => "0101",
		173 => "0101",
		174 => "0101",
		175 => "0101",
		176 => "0100",
		177 => "0100",
		178 => "0100",
		179 => "0100",
		180 => "0100",
		181 => "0100",
		182 => "0100",
		183 => "0100",
		184 => "0100",
		185 => "0100",
		186 => "0100",
		187 => "0100",
		188 => "0100",
		189 => "0100",
		190 => "0100",
		191 => "0100",
		192 => "0011",
		193 => "0011",
		194 => "0011",
		195 => "0011",
		196 => "0011",
		197 => "0011",
		198 => "0011",
		199 => "0011",
		200 => "0011",
		201 => "0011",
		202 => "0011",
		203 => "0011",
		204 => "0011",
		205 => "0011",
		206 => "0011",
		207 => "0011",
		208 => "0010",
		209 => "0010",
		210 => "0010",
		211 => "0010",
		212 => "0010",
		213 => "0010",
		214 => "0010",
		215 => "0010",
		216 => "0010",
		217 => "0010",
		218 => "0010",
		219 => "0010",
		220 => "0010",
		221 => "0010",
		222 => "0010",
		223 => "0010",
		224 => "0001",
		225 => "0001",
		226 => "0001",
		227 => "0001",
		228 => "0001",
		229 => "0001",
		230 => "0001",
		231 => "0001",
		232 => "0001",
		233 => "0001",
		234 => "0001",
		235 => "0001",
		236 => "0001",
		237 => "0001",
		238 => "0001",
		239 => "0001",
		240 => "0000",
		241 => "0000",
		242 => "0000",
		243 => "0000",
		244 => "0000",
		245 => "0000",
		246 => "0000",
		247 => "0000",
		248 => "0000",
		249 => "0000",
		250 => "0000",
		251 => "0000",
		252 => "0000",
		253 => "0000",
		254 => "0000",
		255 => "0000"
	);

begin

	value <= ROM( to_integer( unsigned(address) ) );

end architecture;
